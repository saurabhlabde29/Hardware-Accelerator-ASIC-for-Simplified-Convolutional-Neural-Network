
module macopertion_1_DW02_mac_1 ( A, B, C, TC, MAC );
  input [15:0] A;
  input [15:0] B;
  input [31:0] C;
  output [31:0] MAC;
  input TC;
  wire   n6, n12, n18, n24, n30, n36, n42, n48, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n88, n90, n91, n92, n93, n94, n96, n98, n99, n100, n101, n102,
         n104, n106, n107, n108, n109, n110, n112, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n131, n133, n134, n135, n136, n137, n138, n139, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n159, n161, n162, n163, n164, n166, n168,
         n169, n171, n173, n174, n175, n177, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n189, n191, n192, n194, n195, n197, n199,
         n201, n203, n204, n205, n207, n208, n209, n210, n211, n216, n217,
         n221, n222, n223, n224, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n494, n497, n500, n503, n506, n509, n512, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n811, n812, n813, n814, n815, n816, n817, n818, n834, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985;

  FA_X1 U53 ( .A(n223), .B(n222), .CI(n78), .CO(n77), .S(MAC[30]) );
  FA_X1 U54 ( .A(n224), .B(n227), .CI(n79), .CO(n78), .S(MAC[29]) );
  FA_X1 U55 ( .A(n231), .B(n228), .CI(n80), .CO(n79), .S(MAC[28]) );
  FA_X1 U56 ( .A(n237), .B(n232), .CI(n81), .CO(n80), .S(MAC[27]) );
  FA_X1 U58 ( .A(n244), .B(n251), .CI(n83), .CO(n82), .S(MAC[25]) );
  XOR2_X2 U59 ( .A(n52), .B(n86), .Z(MAC[24]) );
  NAND2_X2 U61 ( .A1(n195), .A2(n85), .ZN(n52) );
  NAND2_X2 U64 ( .A1(n252), .A2(n259), .ZN(n85) );
  XNOR2_X2 U65 ( .A(n91), .B(n53), .ZN(MAC[23]) );
  NAND2_X2 U69 ( .A1(n959), .A2(n90), .ZN(n53) );
  NAND2_X2 U72 ( .A1(n260), .A2(n269), .ZN(n90) );
  XOR2_X2 U73 ( .A(n54), .B(n94), .Z(MAC[22]) );
  NAND2_X2 U75 ( .A1(n197), .A2(n93), .ZN(n54) );
  NAND2_X2 U78 ( .A1(n270), .A2(n279), .ZN(n93) );
  XNOR2_X2 U79 ( .A(n99), .B(n55), .ZN(MAC[21]) );
  NAND2_X2 U83 ( .A1(n958), .A2(n98), .ZN(n55) );
  NAND2_X2 U86 ( .A1(n280), .A2(n291), .ZN(n98) );
  XOR2_X2 U87 ( .A(n56), .B(n102), .Z(MAC[20]) );
  NAND2_X2 U89 ( .A1(n199), .A2(n101), .ZN(n56) );
  NAND2_X2 U92 ( .A1(n292), .A2(n303), .ZN(n101) );
  XNOR2_X2 U93 ( .A(n107), .B(n57), .ZN(MAC[19]) );
  NAND2_X2 U97 ( .A1(n957), .A2(n106), .ZN(n57) );
  NAND2_X2 U100 ( .A1(n304), .A2(n317), .ZN(n106) );
  XOR2_X2 U101 ( .A(n58), .B(n110), .Z(MAC[18]) );
  NAND2_X2 U103 ( .A1(n201), .A2(n109), .ZN(n58) );
  NAND2_X2 U106 ( .A1(n318), .A2(n331), .ZN(n109) );
  XNOR2_X2 U107 ( .A(n115), .B(n59), .ZN(MAC[17]) );
  NAND2_X2 U111 ( .A1(n956), .A2(n114), .ZN(n59) );
  NAND2_X2 U114 ( .A1(n332), .A2(n347), .ZN(n114) );
  XOR2_X2 U115 ( .A(n60), .B(n118), .Z(MAC[16]) );
  NAND2_X2 U117 ( .A1(n203), .A2(n117), .ZN(n60) );
  NAND2_X2 U120 ( .A1(n348), .A2(n363), .ZN(n117) );
  XNOR2_X2 U121 ( .A(n123), .B(n61), .ZN(MAC[15]) );
  NAND2_X2 U128 ( .A1(n364), .A2(n379), .ZN(n122) );
  XOR2_X2 U129 ( .A(n62), .B(n126), .Z(MAC[14]) );
  NAND2_X2 U131 ( .A1(n205), .A2(n125), .ZN(n62) );
  NAND2_X2 U134 ( .A1(n380), .A2(n393), .ZN(n125) );
  XOR2_X2 U135 ( .A(n63), .B(n134), .Z(MAC[13]) );
  NAND2_X2 U138 ( .A1(n955), .A2(n135), .ZN(n128) );
  NAND2_X2 U145 ( .A1(n394), .A2(n407), .ZN(n133) );
  XOR2_X2 U146 ( .A(n64), .B(n139), .Z(MAC[12]) );
  NAND2_X2 U150 ( .A1(n207), .A2(n138), .ZN(n64) );
  NAND2_X2 U153 ( .A1(n408), .A2(n419), .ZN(n138) );
  XNOR2_X2 U154 ( .A(n144), .B(n65), .ZN(MAC[11]) );
  NAND2_X2 U161 ( .A1(n420), .A2(n431), .ZN(n143) );
  XNOR2_X2 U162 ( .A(n150), .B(n66), .ZN(MAC[10]) );
  NAND2_X2 U167 ( .A1(n209), .A2(n149), .ZN(n66) );
  XOR2_X2 U171 ( .A(n67), .B(n153), .Z(MAC[9]) );
  NAND2_X2 U173 ( .A1(n210), .A2(n152), .ZN(n67) );
  NAND2_X2 U176 ( .A1(n442), .A2(n451), .ZN(n152) );
  XOR2_X2 U177 ( .A(n157), .B(n68), .Z(MAC[8]) );
  NAND2_X2 U180 ( .A1(n211), .A2(n156), .ZN(n68) );
  NAND2_X2 U183 ( .A1(n452), .A2(n459), .ZN(n156) );
  XNOR2_X2 U184 ( .A(n69), .B(n162), .ZN(MAC[7]) );
  NAND2_X2 U188 ( .A1(n963), .A2(n161), .ZN(n69) );
  NAND2_X2 U191 ( .A1(n460), .A2(n467), .ZN(n161) );
  XOR2_X2 U192 ( .A(n70), .B(n169), .Z(MAC[6]) );
  NAND2_X2 U194 ( .A1(n961), .A2(n962), .ZN(n163) );
  NAND2_X2 U198 ( .A1(n961), .A2(n168), .ZN(n70) );
  NAND2_X2 U201 ( .A1(n468), .A2(n473), .ZN(n168) );
  XNOR2_X2 U202 ( .A(n174), .B(n71), .ZN(MAC[5]) );
  NAND2_X2 U206 ( .A1(n962), .A2(n173), .ZN(n71) );
  NAND2_X2 U209 ( .A1(n474), .A2(n479), .ZN(n173) );
  XNOR2_X2 U210 ( .A(n72), .B(n180), .ZN(MAC[4]) );
  NAND2_X2 U215 ( .A1(n960), .A2(n179), .ZN(n72) );
  NAND2_X2 U218 ( .A1(n480), .A2(n483), .ZN(n179) );
  XOR2_X2 U219 ( .A(n183), .B(n73), .Z(MAC[3]) );
  NAND2_X2 U221 ( .A1(n216), .A2(n182), .ZN(n73) );
  NAND2_X2 U224 ( .A1(n484), .A2(n486), .ZN(n182) );
  XOR2_X2 U225 ( .A(n187), .B(n74), .Z(MAC[2]) );
  NAND2_X2 U228 ( .A1(n217), .A2(n186), .ZN(n74) );
  NAND2_X2 U231 ( .A1(n488), .A2(n489), .ZN(n186) );
  XNOR2_X2 U232 ( .A(n75), .B(n192), .ZN(MAC[1]) );
  NAND2_X2 U236 ( .A1(n964), .A2(n191), .ZN(n75) );
  NAND2_X2 U239 ( .A1(n490), .A2(n522), .ZN(n191) );
  NAND2_X2 U245 ( .A1(n658), .A2(C[0]), .ZN(n194) );
  FA_X1 U247 ( .A(C[29]), .B(C[30]), .CI(n523), .CO(n221), .S(n222) );
  FA_X1 U248 ( .A(n524), .B(n226), .CI(n229), .CO(n223), .S(n224) );
  FA_X1 U250 ( .A(n233), .B(n540), .CI(n230), .CO(n227), .S(n228) );
  FA_X1 U251 ( .A(C[27]), .B(C[28]), .CI(n525), .CO(n229), .S(n230) );
  FA_X1 U252 ( .A(n234), .B(n241), .CI(n239), .CO(n231), .S(n232) );
  FA_X1 U253 ( .A(n541), .B(n236), .CI(n526), .CO(n233), .S(n234) );
  FA_X1 U255 ( .A(n245), .B(n242), .CI(n240), .CO(n237), .S(n238) );
  FA_X1 U256 ( .A(n557), .B(n527), .CI(n247), .CO(n239), .S(n240) );
  FA_X1 U257 ( .A(C[25]), .B(C[26]), .CI(n542), .CO(n241), .S(n242) );
  FA_X1 U258 ( .A(n246), .B(n248), .CI(n253), .CO(n243), .S(n244) );
  FA_X1 U259 ( .A(n257), .B(n528), .CI(n255), .CO(n245), .S(n246) );
  FA_X1 U260 ( .A(n558), .B(n250), .CI(n543), .CO(n247), .S(n248) );
  FA_X1 U262 ( .A(n254), .B(n263), .CI(n261), .CO(n251), .S(n252) );
  FA_X1 U263 ( .A(n258), .B(n265), .CI(n256), .CO(n253), .S(n254) );
  FA_X1 U264 ( .A(n544), .B(n529), .CI(n574), .CO(n255), .S(n256) );
  FA_X1 U265 ( .A(C[23]), .B(C[24]), .CI(n559), .CO(n257), .S(n258) );
  FA_X1 U266 ( .A(n271), .B(n264), .CI(n262), .CO(n259), .S(n260) );
  FA_X1 U267 ( .A(n266), .B(n275), .CI(n273), .CO(n261), .S(n262) );
  FA_X1 U268 ( .A(n530), .B(n545), .CI(n277), .CO(n263), .S(n264) );
  FA_X1 U269 ( .A(n575), .B(n268), .CI(n560), .CO(n265), .S(n266) );
  FA_X1 U271 ( .A(n281), .B(n274), .CI(n272), .CO(n269), .S(n270) );
  FA_X1 U272 ( .A(n276), .B(n278), .CI(n283), .CO(n271), .S(n272) );
  FA_X1 U273 ( .A(n287), .B(n576), .CI(n285), .CO(n273), .S(n274) );
  FA_X1 U274 ( .A(n531), .B(n546), .CI(n591), .CO(n275), .S(n276) );
  FA_X1 U275 ( .A(C[21]), .B(C[22]), .CI(n561), .CO(n277), .S(n278) );
  FA_X1 U276 ( .A(n293), .B(n284), .CI(n282), .CO(n279), .S(n280) );
  FA_X1 U277 ( .A(n297), .B(n286), .CI(n295), .CO(n281), .S(n282) );
  FA_X1 U278 ( .A(n299), .B(n301), .CI(n288), .CO(n283), .S(n284) );
  FA_X1 U279 ( .A(n547), .B(n532), .CI(n562), .CO(n285), .S(n286) );
  FA_X1 U280 ( .A(n592), .B(n290), .CI(n577), .CO(n287), .S(n288) );
  FA_X1 U282 ( .A(n305), .B(n296), .CI(n294), .CO(n291), .S(n292) );
  FA_X1 U283 ( .A(n298), .B(n309), .CI(n307), .CO(n293), .S(n294) );
  FA_X1 U284 ( .A(n302), .B(n311), .CI(n300), .CO(n295), .S(n296) );
  FA_X1 U285 ( .A(n533), .B(n548), .CI(n313), .CO(n297), .S(n298) );
  FA_X1 U286 ( .A(n593), .B(n563), .CI(n608), .CO(n299), .S(n300) );
  FA_X1 U287 ( .A(C[19]), .B(C[20]), .CI(n578), .CO(n301), .S(n302) );
  FA_X1 U288 ( .A(n319), .B(n308), .CI(n306), .CO(n303), .S(n304) );
  FA_X1 U289 ( .A(n310), .B(n323), .CI(n321), .CO(n305), .S(n306) );
  FA_X1 U290 ( .A(n314), .B(n325), .CI(n312), .CO(n307), .S(n308) );
  FA_X1 U291 ( .A(n329), .B(n549), .CI(n327), .CO(n309), .S(n310) );
  FA_X1 U292 ( .A(n534), .B(n579), .CI(n564), .CO(n311), .S(n312) );
  FA_X1 U293 ( .A(n609), .B(n316), .CI(n594), .CO(n313), .S(n314) );
  FA_X1 U295 ( .A(n333), .B(n322), .CI(n320), .CO(n317), .S(n318) );
  FA_X1 U296 ( .A(n324), .B(n337), .CI(n335), .CO(n319), .S(n320) );
  FA_X1 U297 ( .A(n326), .B(n330), .CI(n328), .CO(n321), .S(n322) );
  FA_X1 U298 ( .A(n341), .B(n343), .CI(n339), .CO(n323), .S(n324) );
  FA_X1 U299 ( .A(n550), .B(n610), .CI(n595), .CO(n325), .S(n326) );
  FA_X1 U300 ( .A(n535), .B(n565), .CI(n625), .CO(n327), .S(n328) );
  FA_X1 U301 ( .A(C[17]), .B(C[18]), .CI(n580), .CO(n329), .S(n330) );
  FA_X1 U302 ( .A(n349), .B(n336), .CI(n334), .CO(n331), .S(n332) );
  FA_X1 U303 ( .A(n338), .B(n353), .CI(n351), .CO(n333), .S(n334) );
  FA_X1 U304 ( .A(n342), .B(n344), .CI(n340), .CO(n335), .S(n336) );
  FA_X1 U305 ( .A(n357), .B(n359), .CI(n355), .CO(n337), .S(n338) );
  FA_X1 U306 ( .A(n566), .B(n581), .CI(n361), .CO(n339), .S(n340) );
  FA_X1 U307 ( .A(n536), .B(n596), .CI(n551), .CO(n341), .S(n342) );
  FA_X1 U308 ( .A(n626), .B(n346), .CI(n611), .CO(n343), .S(n344) );
  FA_X1 U310 ( .A(n365), .B(n352), .CI(n350), .CO(n347), .S(n348) );
  FA_X1 U311 ( .A(n354), .B(n369), .CI(n367), .CO(n349), .S(n350) );
  FA_X1 U312 ( .A(n371), .B(n360), .CI(n356), .CO(n351), .S(n352) );
  FA_X1 U313 ( .A(n373), .B(n375), .CI(n358), .CO(n353), .S(n354) );
  FA_X1 U314 ( .A(n377), .B(n582), .CI(n362), .CO(n355), .S(n356) );
  FA_X1 U315 ( .A(n537), .B(n612), .CI(n552), .CO(n357), .S(n358) );
  FA_X1 U316 ( .A(n627), .B(n567), .CI(n642), .CO(n359), .S(n360) );
  XNOR2_X2 U317 ( .A(n597), .B(C[16]), .ZN(n362) );
  OR2_X2 U318 ( .A1(n597), .A2(C[16]), .ZN(n361) );
  FA_X1 U319 ( .A(n381), .B(n368), .CI(n366), .CO(n363), .S(n364) );
  FA_X1 U320 ( .A(n383), .B(n372), .CI(n370), .CO(n365), .S(n366) );
  FA_X1 U321 ( .A(n376), .B(n374), .CI(n385), .CO(n367), .S(n368) );
  FA_X1 U322 ( .A(n389), .B(n378), .CI(n387), .CO(n369), .S(n370) );
  FA_X1 U323 ( .A(n598), .B(n613), .CI(n391), .CO(n371), .S(n372) );
  FA_X1 U324 ( .A(n553), .B(n568), .CI(n583), .CO(n373), .S(n374) );
  FA_X1 U325 ( .A(n515), .B(n643), .CI(n628), .CO(n375), .S(n376) );
  HA_X1 U326 ( .A(C[15]), .B(n538), .CO(n377), .S(n378) );
  FA_X1 U327 ( .A(n395), .B(n384), .CI(n382), .CO(n379), .S(n380) );
  FA_X1 U328 ( .A(n397), .B(n399), .CI(n386), .CO(n381), .S(n382) );
  FA_X1 U330 ( .A(n403), .B(n405), .CI(n401), .CO(n385), .S(n386) );
  FA_X1 U331 ( .A(n584), .B(n614), .CI(n599), .CO(n387), .S(n388) );
  FA_X1 U332 ( .A(n554), .B(n629), .CI(n569), .CO(n389), .S(n390) );
  FA_X1 U333 ( .A(n539), .B(C[14]), .CI(n644), .CO(n391), .S(n392) );
  FA_X1 U334 ( .A(n398), .B(n409), .CI(n396), .CO(n393), .S(n394) );
  FA_X1 U335 ( .A(n411), .B(n404), .CI(n400), .CO(n395), .S(n396) );
  FA_X1 U336 ( .A(n413), .B(n415), .CI(n402), .CO(n397), .S(n398) );
  FA_X1 U337 ( .A(n417), .B(n615), .CI(n406), .CO(n399), .S(n400) );
  FA_X1 U338 ( .A(n630), .B(n585), .CI(n600), .CO(n401), .S(n402) );
  FA_X1 U339 ( .A(n516), .B(n645), .CI(n570), .CO(n403), .S(n404) );
  HA_X1 U340 ( .A(C[13]), .B(n555), .CO(n405), .S(n406) );
  FA_X1 U341 ( .A(n421), .B(n412), .CI(n410), .CO(n407), .S(n408) );
  FA_X1 U342 ( .A(n414), .B(n416), .CI(n423), .CO(n409), .S(n410) );
  FA_X1 U343 ( .A(n425), .B(n427), .CI(n418), .CO(n411), .S(n412) );
  FA_X1 U344 ( .A(n601), .B(n616), .CI(n429), .CO(n413), .S(n414) );
  FA_X1 U345 ( .A(n571), .B(n631), .CI(n586), .CO(n415), .S(n416) );
  FA_X1 U346 ( .A(n556), .B(C[12]), .CI(n646), .CO(n417), .S(n418) );
  FA_X1 U347 ( .A(n433), .B(n424), .CI(n422), .CO(n419), .S(n420) );
  FA_X1 U348 ( .A(n428), .B(n426), .CI(n435), .CO(n421), .S(n422) );
  FA_X1 U349 ( .A(n430), .B(n439), .CI(n437), .CO(n423), .S(n424) );
  FA_X1 U350 ( .A(n587), .B(n617), .CI(n602), .CO(n425), .S(n426) );
  FA_X1 U351 ( .A(n517), .B(n647), .CI(n632), .CO(n427), .S(n428) );
  HA_X1 U352 ( .A(C[11]), .B(n572), .CO(n429), .S(n430) );
  FA_X1 U353 ( .A(n443), .B(n436), .CI(n434), .CO(n431), .S(n432) );
  FA_X1 U354 ( .A(n438), .B(n440), .CI(n445), .CO(n433), .S(n434) );
  FA_X1 U355 ( .A(n449), .B(n618), .CI(n447), .CO(n435), .S(n436) );
  FA_X1 U356 ( .A(n588), .B(n633), .CI(n603), .CO(n437), .S(n438) );
  FA_X1 U357 ( .A(n573), .B(C[10]), .CI(n648), .CO(n439), .S(n440) );
  FA_X1 U358 ( .A(n453), .B(n446), .CI(n444), .CO(n441), .S(n442) );
  FA_X1 U359 ( .A(n455), .B(n450), .CI(n448), .CO(n443), .S(n444) );
  FA_X1 U360 ( .A(n604), .B(n619), .CI(n457), .CO(n445), .S(n446) );
  FA_X1 U361 ( .A(n518), .B(n649), .CI(n634), .CO(n447), .S(n448) );
  HA_X1 U362 ( .A(C[9]), .B(n589), .CO(n449), .S(n450) );
  FA_X1 U363 ( .A(n461), .B(n456), .CI(n454), .CO(n451), .S(n452) );
  FA_X1 U364 ( .A(n463), .B(n465), .CI(n458), .CO(n453), .S(n454) );
  FA_X1 U365 ( .A(n605), .B(n635), .CI(n620), .CO(n455), .S(n456) );
  FA_X1 U366 ( .A(n590), .B(C[8]), .CI(n650), .CO(n457), .S(n458) );
  FA_X1 U367 ( .A(n464), .B(n469), .CI(n462), .CO(n459), .S(n460) );
  FA_X1 U368 ( .A(n471), .B(n636), .CI(n466), .CO(n461), .S(n462) );
  FA_X1 U369 ( .A(n519), .B(n651), .CI(n621), .CO(n463), .S(n464) );
  HA_X1 U370 ( .A(C[7]), .B(n606), .CO(n465), .S(n466) );
  FA_X1 U371 ( .A(n472), .B(n475), .CI(n470), .CO(n467), .S(n468) );
  FA_X1 U372 ( .A(n622), .B(n637), .CI(n477), .CO(n469), .S(n470) );
  FA_X1 U373 ( .A(n607), .B(C[6]), .CI(n652), .CO(n471), .S(n472) );
  FA_X1 U374 ( .A(n478), .B(n481), .CI(n476), .CO(n473), .S(n474) );
  FA_X1 U375 ( .A(n520), .B(n653), .CI(n638), .CO(n475), .S(n476) );
  HA_X1 U376 ( .A(C[5]), .B(n623), .CO(n477), .S(n478) );
  FA_X1 U377 ( .A(n485), .B(n639), .CI(n482), .CO(n479), .S(n480) );
  FA_X1 U378 ( .A(n624), .B(C[4]), .CI(n654), .CO(n481), .S(n482) );
  FA_X1 U379 ( .A(n521), .B(n640), .CI(n487), .CO(n483), .S(n484) );
  HA_X1 U380 ( .A(C[3]), .B(n655), .CO(n485), .S(n486) );
  FA_X1 U381 ( .A(n641), .B(C[2]), .CI(n656), .CO(n487), .S(n488) );
  HA_X1 U382 ( .A(C[1]), .B(n657), .CO(n489), .S(n490) );
  OAI22_X2 U383 ( .A1(n48), .A2(n985), .B1(n675), .B2(n971), .ZN(n515) );
  OAI22_X2 U386 ( .A1(n48), .A2(n660), .B1(n971), .B2(n659), .ZN(n524) );
  OAI22_X2 U387 ( .A1(n48), .A2(n661), .B1(n971), .B2(n660), .ZN(n525) );
  OAI22_X2 U388 ( .A1(n48), .A2(n662), .B1(n971), .B2(n661), .ZN(n526) );
  OAI22_X2 U389 ( .A1(n48), .A2(n663), .B1(n971), .B2(n662), .ZN(n527) );
  OAI22_X2 U390 ( .A1(n48), .A2(n664), .B1(n971), .B2(n663), .ZN(n528) );
  OAI22_X2 U392 ( .A1(n48), .A2(n666), .B1(n971), .B2(n665), .ZN(n530) );
  OAI22_X2 U393 ( .A1(n48), .A2(n667), .B1(n971), .B2(n666), .ZN(n531) );
  OAI22_X2 U394 ( .A1(n48), .A2(n668), .B1(n971), .B2(n667), .ZN(n532) );
  OAI22_X2 U395 ( .A1(n48), .A2(n669), .B1(n971), .B2(n668), .ZN(n533) );
  OAI22_X2 U396 ( .A1(n48), .A2(n670), .B1(n971), .B2(n669), .ZN(n534) );
  OAI22_X2 U397 ( .A1(n48), .A2(n671), .B1(n971), .B2(n670), .ZN(n535) );
  OAI22_X2 U398 ( .A1(n48), .A2(n672), .B1(n971), .B2(n671), .ZN(n536) );
  OAI22_X2 U399 ( .A1(n48), .A2(n673), .B1(n971), .B2(n672), .ZN(n537) );
  OAI22_X2 U400 ( .A1(n48), .A2(n674), .B1(n971), .B2(n673), .ZN(n538) );
  AND2_X2 U401 ( .A1(B[0]), .A2(n948), .ZN(n539) );
  XNOR2_X2 U403 ( .A(A[15]), .B(B[15]), .ZN(n659) );
  XNOR2_X2 U404 ( .A(A[15]), .B(B[14]), .ZN(n660) );
  XNOR2_X2 U405 ( .A(A[15]), .B(B[13]), .ZN(n661) );
  XNOR2_X2 U406 ( .A(A[15]), .B(B[12]), .ZN(n662) );
  XNOR2_X2 U407 ( .A(A[15]), .B(B[11]), .ZN(n663) );
  XNOR2_X2 U408 ( .A(A[15]), .B(B[10]), .ZN(n664) );
  XNOR2_X2 U409 ( .A(A[15]), .B(B[9]), .ZN(n665) );
  XNOR2_X2 U410 ( .A(A[15]), .B(B[8]), .ZN(n666) );
  XNOR2_X2 U411 ( .A(A[15]), .B(B[7]), .ZN(n667) );
  XNOR2_X2 U412 ( .A(A[15]), .B(B[6]), .ZN(n668) );
  XNOR2_X2 U413 ( .A(A[15]), .B(B[5]), .ZN(n669) );
  XNOR2_X2 U414 ( .A(A[15]), .B(B[4]), .ZN(n670) );
  XNOR2_X2 U416 ( .A(A[15]), .B(B[2]), .ZN(n672) );
  XNOR2_X2 U417 ( .A(A[15]), .B(B[1]), .ZN(n673) );
  XNOR2_X2 U418 ( .A(B[0]), .B(A[15]), .ZN(n674) );
  OR2_X2 U419 ( .A1(B[0]), .A2(n985), .ZN(n675) );
  OAI22_X2 U421 ( .A1(n42), .A2(n984), .B1(n692), .B2(n970), .ZN(n516) );
  OAI22_X2 U424 ( .A1(n42), .A2(n677), .B1(n970), .B2(n676), .ZN(n541) );
  OAI22_X2 U425 ( .A1(n42), .A2(n678), .B1(n970), .B2(n677), .ZN(n542) );
  OAI22_X2 U426 ( .A1(n42), .A2(n679), .B1(n970), .B2(n678), .ZN(n543) );
  OAI22_X2 U427 ( .A1(n42), .A2(n680), .B1(n970), .B2(n679), .ZN(n544) );
  OAI22_X2 U428 ( .A1(n42), .A2(n681), .B1(n970), .B2(n680), .ZN(n545) );
  OAI22_X2 U430 ( .A1(n42), .A2(n683), .B1(n970), .B2(n682), .ZN(n547) );
  OAI22_X2 U431 ( .A1(n42), .A2(n684), .B1(n970), .B2(n683), .ZN(n548) );
  OAI22_X2 U432 ( .A1(n42), .A2(n685), .B1(n970), .B2(n684), .ZN(n549) );
  OAI22_X2 U433 ( .A1(n42), .A2(n686), .B1(n970), .B2(n685), .ZN(n550) );
  OAI22_X2 U434 ( .A1(n42), .A2(n687), .B1(n970), .B2(n686), .ZN(n551) );
  OAI22_X2 U435 ( .A1(n42), .A2(n688), .B1(n970), .B2(n687), .ZN(n552) );
  OAI22_X2 U436 ( .A1(n42), .A2(n689), .B1(n970), .B2(n688), .ZN(n553) );
  OAI22_X2 U437 ( .A1(n42), .A2(n690), .B1(n970), .B2(n689), .ZN(n554) );
  OAI22_X2 U438 ( .A1(n42), .A2(n691), .B1(n970), .B2(n690), .ZN(n555) );
  AND2_X2 U439 ( .A1(B[0]), .A2(n949), .ZN(n556) );
  XNOR2_X2 U441 ( .A(A[13]), .B(B[15]), .ZN(n676) );
  XNOR2_X2 U442 ( .A(A[13]), .B(B[14]), .ZN(n677) );
  XNOR2_X2 U443 ( .A(A[13]), .B(B[13]), .ZN(n678) );
  XNOR2_X2 U444 ( .A(A[13]), .B(B[12]), .ZN(n679) );
  XNOR2_X2 U445 ( .A(A[13]), .B(B[11]), .ZN(n680) );
  XNOR2_X2 U446 ( .A(A[13]), .B(B[10]), .ZN(n681) );
  XNOR2_X2 U447 ( .A(A[13]), .B(B[9]), .ZN(n682) );
  XNOR2_X2 U448 ( .A(A[13]), .B(B[8]), .ZN(n683) );
  XNOR2_X2 U449 ( .A(A[13]), .B(B[7]), .ZN(n684) );
  XNOR2_X2 U450 ( .A(A[13]), .B(B[6]), .ZN(n685) );
  XNOR2_X2 U451 ( .A(A[13]), .B(B[5]), .ZN(n686) );
  XNOR2_X2 U452 ( .A(A[13]), .B(B[4]), .ZN(n687) );
  XNOR2_X2 U454 ( .A(A[13]), .B(B[2]), .ZN(n689) );
  XNOR2_X2 U455 ( .A(A[13]), .B(B[1]), .ZN(n690) );
  XNOR2_X2 U456 ( .A(B[0]), .B(A[13]), .ZN(n691) );
  OR2_X2 U457 ( .A1(B[0]), .A2(n984), .ZN(n692) );
  OAI22_X2 U459 ( .A1(n36), .A2(n982), .B1(n709), .B2(n969), .ZN(n517) );
  OAI22_X2 U462 ( .A1(n36), .A2(n694), .B1(n969), .B2(n693), .ZN(n558) );
  OAI22_X2 U463 ( .A1(n36), .A2(n695), .B1(n969), .B2(n694), .ZN(n559) );
  OAI22_X2 U464 ( .A1(n36), .A2(n696), .B1(n969), .B2(n695), .ZN(n560) );
  OAI22_X2 U465 ( .A1(n36), .A2(n697), .B1(n969), .B2(n696), .ZN(n561) );
  OAI22_X2 U466 ( .A1(n36), .A2(n698), .B1(n969), .B2(n697), .ZN(n562) );
  OAI22_X2 U467 ( .A1(n36), .A2(n699), .B1(n969), .B2(n698), .ZN(n563) );
  OAI22_X2 U468 ( .A1(n36), .A2(n700), .B1(n969), .B2(n699), .ZN(n564) );
  OAI22_X2 U469 ( .A1(n36), .A2(n701), .B1(n969), .B2(n700), .ZN(n565) );
  OAI22_X2 U470 ( .A1(n36), .A2(n702), .B1(n969), .B2(n701), .ZN(n566) );
  OAI22_X2 U471 ( .A1(n36), .A2(n703), .B1(n969), .B2(n702), .ZN(n567) );
  OAI22_X2 U472 ( .A1(n36), .A2(n704), .B1(n969), .B2(n703), .ZN(n568) );
  OAI22_X2 U473 ( .A1(n36), .A2(n705), .B1(n969), .B2(n704), .ZN(n569) );
  OAI22_X2 U474 ( .A1(n36), .A2(n706), .B1(n969), .B2(n705), .ZN(n570) );
  OAI22_X2 U475 ( .A1(n36), .A2(n707), .B1(n969), .B2(n706), .ZN(n571) );
  OAI22_X2 U476 ( .A1(n36), .A2(n708), .B1(n969), .B2(n707), .ZN(n572) );
  AND2_X2 U477 ( .A1(B[0]), .A2(n951), .ZN(n573) );
  XNOR2_X2 U479 ( .A(n983), .B(B[15]), .ZN(n693) );
  XNOR2_X2 U480 ( .A(n983), .B(B[14]), .ZN(n694) );
  XNOR2_X2 U481 ( .A(n983), .B(B[13]), .ZN(n695) );
  XNOR2_X2 U482 ( .A(n983), .B(B[12]), .ZN(n696) );
  XNOR2_X2 U483 ( .A(n983), .B(B[11]), .ZN(n697) );
  XNOR2_X2 U484 ( .A(n983), .B(B[10]), .ZN(n698) );
  XNOR2_X2 U485 ( .A(n983), .B(B[9]), .ZN(n699) );
  XNOR2_X2 U486 ( .A(n983), .B(B[8]), .ZN(n700) );
  XNOR2_X2 U487 ( .A(n983), .B(B[7]), .ZN(n701) );
  XNOR2_X2 U488 ( .A(n983), .B(B[6]), .ZN(n702) );
  XNOR2_X2 U489 ( .A(n983), .B(B[5]), .ZN(n703) );
  XNOR2_X2 U490 ( .A(n983), .B(B[4]), .ZN(n704) );
  XNOR2_X2 U492 ( .A(n983), .B(B[2]), .ZN(n706) );
  XNOR2_X2 U493 ( .A(n983), .B(B[1]), .ZN(n707) );
  XNOR2_X2 U494 ( .A(B[0]), .B(n983), .ZN(n708) );
  OR2_X2 U495 ( .A1(B[0]), .A2(n982), .ZN(n709) );
  OAI22_X2 U497 ( .A1(n30), .A2(n980), .B1(n726), .B2(n968), .ZN(n518) );
  OAI22_X2 U500 ( .A1(n30), .A2(n711), .B1(n968), .B2(n710), .ZN(n575) );
  OAI22_X2 U501 ( .A1(n30), .A2(n712), .B1(n968), .B2(n711), .ZN(n576) );
  OAI22_X2 U502 ( .A1(n30), .A2(n713), .B1(n968), .B2(n712), .ZN(n577) );
  OAI22_X2 U503 ( .A1(n30), .A2(n714), .B1(n968), .B2(n713), .ZN(n578) );
  OAI22_X2 U504 ( .A1(n30), .A2(n715), .B1(n968), .B2(n714), .ZN(n579) );
  OAI22_X2 U505 ( .A1(n30), .A2(n716), .B1(n968), .B2(n715), .ZN(n580) );
  OAI22_X2 U506 ( .A1(n30), .A2(n717), .B1(n968), .B2(n716), .ZN(n581) );
  OAI22_X2 U507 ( .A1(n30), .A2(n718), .B1(n968), .B2(n717), .ZN(n582) );
  OAI22_X2 U508 ( .A1(n30), .A2(n719), .B1(n968), .B2(n718), .ZN(n583) );
  OAI22_X2 U509 ( .A1(n30), .A2(n720), .B1(n968), .B2(n719), .ZN(n584) );
  OAI22_X2 U510 ( .A1(n30), .A2(n721), .B1(n968), .B2(n720), .ZN(n585) );
  OAI22_X2 U511 ( .A1(n30), .A2(n722), .B1(n968), .B2(n721), .ZN(n586) );
  OAI22_X2 U512 ( .A1(n30), .A2(n723), .B1(n968), .B2(n722), .ZN(n587) );
  OAI22_X2 U513 ( .A1(n30), .A2(n724), .B1(n968), .B2(n723), .ZN(n588) );
  OAI22_X2 U514 ( .A1(n30), .A2(n725), .B1(n968), .B2(n724), .ZN(n589) );
  AND2_X2 U515 ( .A1(B[0]), .A2(n950), .ZN(n590) );
  XNOR2_X2 U517 ( .A(n981), .B(B[15]), .ZN(n710) );
  XNOR2_X2 U518 ( .A(n981), .B(B[14]), .ZN(n711) );
  XNOR2_X2 U519 ( .A(n981), .B(B[13]), .ZN(n712) );
  XNOR2_X2 U520 ( .A(n981), .B(B[12]), .ZN(n713) );
  XNOR2_X2 U521 ( .A(n981), .B(B[11]), .ZN(n714) );
  XNOR2_X2 U522 ( .A(n981), .B(B[10]), .ZN(n715) );
  XNOR2_X2 U523 ( .A(n981), .B(B[9]), .ZN(n716) );
  XNOR2_X2 U524 ( .A(n981), .B(B[8]), .ZN(n717) );
  XNOR2_X2 U525 ( .A(n981), .B(B[7]), .ZN(n718) );
  XNOR2_X2 U526 ( .A(n981), .B(B[6]), .ZN(n719) );
  XNOR2_X2 U527 ( .A(n981), .B(B[5]), .ZN(n720) );
  XNOR2_X2 U528 ( .A(n981), .B(B[4]), .ZN(n721) );
  XNOR2_X2 U530 ( .A(n981), .B(B[2]), .ZN(n723) );
  XNOR2_X2 U531 ( .A(n981), .B(B[1]), .ZN(n724) );
  XNOR2_X2 U532 ( .A(B[0]), .B(n981), .ZN(n725) );
  OR2_X2 U533 ( .A1(B[0]), .A2(n980), .ZN(n726) );
  OAI22_X2 U535 ( .A1(n24), .A2(n978), .B1(n743), .B2(n967), .ZN(n519) );
  OAI22_X2 U538 ( .A1(n24), .A2(n728), .B1(n967), .B2(n727), .ZN(n592) );
  OAI22_X2 U539 ( .A1(n24), .A2(n729), .B1(n967), .B2(n728), .ZN(n593) );
  OAI22_X2 U540 ( .A1(n24), .A2(n730), .B1(n967), .B2(n729), .ZN(n594) );
  OAI22_X2 U541 ( .A1(n24), .A2(n731), .B1(n967), .B2(n730), .ZN(n595) );
  OAI22_X2 U542 ( .A1(n24), .A2(n732), .B1(n967), .B2(n731), .ZN(n596) );
  OAI22_X2 U543 ( .A1(n24), .A2(n733), .B1(n967), .B2(n732), .ZN(n597) );
  OAI22_X2 U544 ( .A1(n24), .A2(n734), .B1(n967), .B2(n733), .ZN(n598) );
  OAI22_X2 U545 ( .A1(n24), .A2(n735), .B1(n967), .B2(n734), .ZN(n599) );
  OAI22_X2 U546 ( .A1(n24), .A2(n736), .B1(n967), .B2(n735), .ZN(n600) );
  OAI22_X2 U547 ( .A1(n24), .A2(n737), .B1(n967), .B2(n736), .ZN(n601) );
  OAI22_X2 U548 ( .A1(n24), .A2(n738), .B1(n967), .B2(n737), .ZN(n602) );
  OAI22_X2 U549 ( .A1(n24), .A2(n739), .B1(n967), .B2(n738), .ZN(n603) );
  OAI22_X2 U550 ( .A1(n24), .A2(n740), .B1(n967), .B2(n739), .ZN(n604) );
  OAI22_X2 U551 ( .A1(n24), .A2(n741), .B1(n967), .B2(n740), .ZN(n605) );
  OAI22_X2 U552 ( .A1(n24), .A2(n742), .B1(n967), .B2(n741), .ZN(n606) );
  AND2_X2 U553 ( .A1(B[0]), .A2(n947), .ZN(n607) );
  XNOR2_X2 U555 ( .A(n979), .B(B[15]), .ZN(n727) );
  XNOR2_X2 U556 ( .A(n979), .B(B[14]), .ZN(n728) );
  XNOR2_X2 U557 ( .A(n979), .B(B[13]), .ZN(n729) );
  XNOR2_X2 U558 ( .A(n979), .B(B[12]), .ZN(n730) );
  XNOR2_X2 U559 ( .A(n979), .B(B[11]), .ZN(n731) );
  XNOR2_X2 U560 ( .A(n979), .B(B[10]), .ZN(n732) );
  XNOR2_X2 U561 ( .A(n979), .B(B[9]), .ZN(n733) );
  XNOR2_X2 U563 ( .A(n979), .B(B[7]), .ZN(n735) );
  XNOR2_X2 U564 ( .A(n979), .B(B[6]), .ZN(n736) );
  XNOR2_X2 U566 ( .A(n979), .B(B[4]), .ZN(n738) );
  XNOR2_X2 U568 ( .A(n979), .B(B[2]), .ZN(n740) );
  XNOR2_X2 U569 ( .A(n979), .B(B[1]), .ZN(n741) );
  XNOR2_X2 U570 ( .A(B[0]), .B(n979), .ZN(n742) );
  OR2_X2 U571 ( .A1(B[0]), .A2(n978), .ZN(n743) );
  OAI22_X2 U573 ( .A1(n18), .A2(n976), .B1(n760), .B2(n966), .ZN(n520) );
  OAI22_X2 U576 ( .A1(n18), .A2(n745), .B1(n966), .B2(n744), .ZN(n609) );
  OAI22_X2 U577 ( .A1(n18), .A2(n746), .B1(n966), .B2(n745), .ZN(n610) );
  OAI22_X2 U578 ( .A1(n18), .A2(n747), .B1(n966), .B2(n746), .ZN(n611) );
  OAI22_X2 U579 ( .A1(n18), .A2(n748), .B1(n966), .B2(n747), .ZN(n612) );
  OAI22_X2 U580 ( .A1(n18), .A2(n749), .B1(n966), .B2(n748), .ZN(n613) );
  OAI22_X2 U581 ( .A1(n18), .A2(n750), .B1(n966), .B2(n749), .ZN(n614) );
  OAI22_X2 U582 ( .A1(n18), .A2(n751), .B1(n966), .B2(n750), .ZN(n615) );
  OAI22_X2 U583 ( .A1(n18), .A2(n752), .B1(n966), .B2(n751), .ZN(n616) );
  OAI22_X2 U584 ( .A1(n18), .A2(n753), .B1(n966), .B2(n752), .ZN(n617) );
  OAI22_X2 U585 ( .A1(n18), .A2(n754), .B1(n966), .B2(n753), .ZN(n618) );
  OAI22_X2 U586 ( .A1(n18), .A2(n755), .B1(n966), .B2(n754), .ZN(n619) );
  OAI22_X2 U587 ( .A1(n18), .A2(n756), .B1(n966), .B2(n755), .ZN(n620) );
  OAI22_X2 U588 ( .A1(n18), .A2(n757), .B1(n966), .B2(n756), .ZN(n621) );
  OAI22_X2 U589 ( .A1(n18), .A2(n758), .B1(n966), .B2(n757), .ZN(n622) );
  OAI22_X2 U590 ( .A1(n18), .A2(n759), .B1(n966), .B2(n758), .ZN(n623) );
  AND2_X2 U591 ( .A1(B[0]), .A2(n946), .ZN(n624) );
  XNOR2_X2 U593 ( .A(n977), .B(B[15]), .ZN(n744) );
  XNOR2_X2 U594 ( .A(n977), .B(B[14]), .ZN(n745) );
  XNOR2_X2 U595 ( .A(n977), .B(B[13]), .ZN(n746) );
  XNOR2_X2 U596 ( .A(n977), .B(B[12]), .ZN(n747) );
  XNOR2_X2 U597 ( .A(n977), .B(B[11]), .ZN(n748) );
  XNOR2_X2 U598 ( .A(n977), .B(B[10]), .ZN(n749) );
  XNOR2_X2 U599 ( .A(n977), .B(B[9]), .ZN(n750) );
  XNOR2_X2 U600 ( .A(n977), .B(B[8]), .ZN(n751) );
  XNOR2_X2 U601 ( .A(n977), .B(B[7]), .ZN(n752) );
  XNOR2_X2 U602 ( .A(n977), .B(B[6]), .ZN(n753) );
  XNOR2_X2 U603 ( .A(n977), .B(B[5]), .ZN(n754) );
  XNOR2_X2 U604 ( .A(n977), .B(B[4]), .ZN(n755) );
  XNOR2_X2 U606 ( .A(n977), .B(B[2]), .ZN(n757) );
  XNOR2_X2 U607 ( .A(n977), .B(B[1]), .ZN(n758) );
  XNOR2_X2 U608 ( .A(B[0]), .B(n977), .ZN(n759) );
  OR2_X2 U609 ( .A1(B[0]), .A2(n976), .ZN(n760) );
  OAI22_X2 U614 ( .A1(n12), .A2(n762), .B1(n965), .B2(n761), .ZN(n626) );
  OAI22_X2 U615 ( .A1(n12), .A2(n763), .B1(n965), .B2(n762), .ZN(n627) );
  OAI22_X2 U616 ( .A1(n12), .A2(n764), .B1(n965), .B2(n763), .ZN(n628) );
  OAI22_X2 U617 ( .A1(n12), .A2(n765), .B1(n965), .B2(n764), .ZN(n629) );
  OAI22_X2 U618 ( .A1(n12), .A2(n766), .B1(n965), .B2(n765), .ZN(n630) );
  OAI22_X2 U619 ( .A1(n12), .A2(n767), .B1(n965), .B2(n766), .ZN(n631) );
  OAI22_X2 U620 ( .A1(n12), .A2(n768), .B1(n965), .B2(n767), .ZN(n632) );
  OAI22_X2 U621 ( .A1(n12), .A2(n769), .B1(n965), .B2(n768), .ZN(n633) );
  OAI22_X2 U622 ( .A1(n12), .A2(n770), .B1(n965), .B2(n769), .ZN(n634) );
  OAI22_X2 U623 ( .A1(n12), .A2(n771), .B1(n965), .B2(n770), .ZN(n635) );
  OAI22_X2 U624 ( .A1(n12), .A2(n772), .B1(n965), .B2(n771), .ZN(n636) );
  OAI22_X2 U625 ( .A1(n12), .A2(n773), .B1(n965), .B2(n772), .ZN(n637) );
  OAI22_X2 U626 ( .A1(n12), .A2(n774), .B1(n965), .B2(n773), .ZN(n638) );
  OAI22_X2 U627 ( .A1(n12), .A2(n775), .B1(n965), .B2(n774), .ZN(n639) );
  OAI22_X2 U628 ( .A1(n12), .A2(n776), .B1(n965), .B2(n775), .ZN(n640) );
  AND2_X2 U629 ( .A1(B[0]), .A2(n945), .ZN(n641) );
  XNOR2_X2 U631 ( .A(n975), .B(B[15]), .ZN(n761) );
  XNOR2_X2 U632 ( .A(n975), .B(B[14]), .ZN(n762) );
  XNOR2_X2 U633 ( .A(n975), .B(B[13]), .ZN(n763) );
  XNOR2_X2 U634 ( .A(n975), .B(B[12]), .ZN(n764) );
  XNOR2_X2 U635 ( .A(n975), .B(B[11]), .ZN(n765) );
  XNOR2_X2 U636 ( .A(n975), .B(B[10]), .ZN(n766) );
  XNOR2_X2 U637 ( .A(n975), .B(B[9]), .ZN(n767) );
  XNOR2_X2 U639 ( .A(n975), .B(B[7]), .ZN(n769) );
  XNOR2_X2 U640 ( .A(n975), .B(B[6]), .ZN(n770) );
  XNOR2_X2 U642 ( .A(n975), .B(B[4]), .ZN(n772) );
  XNOR2_X2 U644 ( .A(n975), .B(B[2]), .ZN(n774) );
  XNOR2_X2 U645 ( .A(n975), .B(B[1]), .ZN(n775) );
  XNOR2_X2 U646 ( .A(B[0]), .B(n975), .ZN(n776) );
  OR2_X2 U647 ( .A1(B[0]), .A2(n974), .ZN(n777) );
  OAI22_X2 U649 ( .A1(n6), .A2(n972), .B1(n794), .B2(n834), .ZN(n522) );
  OAI22_X2 U652 ( .A1(n6), .A2(n779), .B1(n778), .B2(n834), .ZN(n643) );
  OAI22_X2 U653 ( .A1(n6), .A2(n780), .B1(n779), .B2(n834), .ZN(n644) );
  OAI22_X2 U654 ( .A1(n6), .A2(n781), .B1(n780), .B2(n834), .ZN(n645) );
  OAI22_X2 U655 ( .A1(n6), .A2(n782), .B1(n781), .B2(n834), .ZN(n646) );
  OAI22_X2 U656 ( .A1(n6), .A2(n783), .B1(n782), .B2(n834), .ZN(n647) );
  OAI22_X2 U657 ( .A1(n6), .A2(n784), .B1(n783), .B2(n834), .ZN(n648) );
  OAI22_X2 U658 ( .A1(n6), .A2(n785), .B1(n784), .B2(n834), .ZN(n649) );
  OAI22_X2 U659 ( .A1(n6), .A2(n786), .B1(n785), .B2(n834), .ZN(n650) );
  OAI22_X2 U660 ( .A1(n6), .A2(n787), .B1(n786), .B2(n834), .ZN(n651) );
  OAI22_X2 U661 ( .A1(n6), .A2(n788), .B1(n787), .B2(n834), .ZN(n652) );
  OAI22_X2 U662 ( .A1(n6), .A2(n789), .B1(n788), .B2(n834), .ZN(n653) );
  OAI22_X2 U663 ( .A1(n6), .A2(n790), .B1(n789), .B2(n834), .ZN(n654) );
  OAI22_X2 U665 ( .A1(n6), .A2(n792), .B1(n791), .B2(n834), .ZN(n656) );
  OAI22_X2 U666 ( .A1(n6), .A2(n793), .B1(n792), .B2(n834), .ZN(n657) );
  AND2_X2 U667 ( .A1(B[0]), .A2(A[0]), .ZN(n658) );
  XNOR2_X2 U669 ( .A(n973), .B(B[15]), .ZN(n778) );
  XNOR2_X2 U670 ( .A(n973), .B(B[14]), .ZN(n779) );
  XNOR2_X2 U671 ( .A(n973), .B(B[13]), .ZN(n780) );
  XNOR2_X2 U672 ( .A(n973), .B(B[12]), .ZN(n781) );
  XNOR2_X2 U673 ( .A(n973), .B(B[11]), .ZN(n782) );
  XNOR2_X2 U674 ( .A(n973), .B(B[10]), .ZN(n783) );
  XNOR2_X2 U675 ( .A(n973), .B(B[9]), .ZN(n784) );
  XNOR2_X2 U677 ( .A(n973), .B(B[7]), .ZN(n786) );
  XNOR2_X2 U678 ( .A(n973), .B(B[6]), .ZN(n787) );
  XNOR2_X2 U680 ( .A(n973), .B(B[4]), .ZN(n789) );
  XNOR2_X2 U682 ( .A(n973), .B(B[2]), .ZN(n791) );
  XNOR2_X2 U683 ( .A(n973), .B(B[1]), .ZN(n792) );
  XNOR2_X2 U684 ( .A(B[0]), .B(n973), .ZN(n793) );
  OR2_X2 U685 ( .A1(B[0]), .A2(n972), .ZN(n794) );
  XOR2_X2 U711 ( .A(A[14]), .B(A[15]), .Z(n811) );
  XOR2_X2 U714 ( .A(A[12]), .B(A[13]), .Z(n812) );
  XOR2_X2 U717 ( .A(A[10]), .B(n983), .Z(n813) );
  XOR2_X2 U720 ( .A(A[8]), .B(n981), .Z(n814) );
  XOR2_X2 U723 ( .A(A[6]), .B(n979), .Z(n815) );
  XOR2_X2 U726 ( .A(A[4]), .B(n977), .Z(n816) );
  XOR2_X2 U729 ( .A(A[2]), .B(n975), .Z(n817) );
  XOR2_X2 U732 ( .A(A[0]), .B(n973), .Z(n818) );
  AOI21_X2 U737 ( .B1(n127), .B2(n119), .A(n120), .ZN(n118) );
  XOR2_X2 U738 ( .A(n238), .B(n243), .Z(n937) );
  XOR2_X2 U739 ( .A(n82), .B(n937), .Z(MAC[26]) );
  NAND2_X2 U740 ( .A1(n238), .A2(n82), .ZN(n938) );
  NAND2_X2 U741 ( .A1(n243), .A2(n82), .ZN(n939) );
  NAND2_X2 U742 ( .A1(n243), .A2(n238), .ZN(n940) );
  NAND3_X2 U743 ( .A1(n940), .A2(n939), .A3(n938), .ZN(n81) );
  XOR2_X2 U744 ( .A(n390), .B(n392), .Z(n941) );
  XOR2_X2 U745 ( .A(n388), .B(n941), .Z(n384) );
  NAND2_X2 U746 ( .A1(n390), .A2(n388), .ZN(n942) );
  NAND2_X2 U747 ( .A1(n392), .A2(n388), .ZN(n943) );
  NAND2_X2 U748 ( .A1(n392), .A2(n390), .ZN(n944) );
  NAND3_X2 U749 ( .A1(n944), .A2(n943), .A3(n942), .ZN(n383) );
  XNOR2_X1 U750 ( .A(n975), .B(B[8]), .ZN(n768) );
  XNOR2_X1 U751 ( .A(n975), .B(B[5]), .ZN(n771) );
  XNOR2_X1 U752 ( .A(n973), .B(B[5]), .ZN(n788) );
  XNOR2_X1 U753 ( .A(n973), .B(B[8]), .ZN(n785) );
  XNOR2_X1 U754 ( .A(n979), .B(B[8]), .ZN(n734) );
  XNOR2_X1 U755 ( .A(n979), .B(B[5]), .ZN(n737) );
  OAI22_X1 U756 ( .A1(n12), .A2(n974), .B1(n777), .B2(n965), .ZN(n521) );
  INV_X1 U757 ( .A(A[13]), .ZN(n984) );
  XOR2_X2 U758 ( .A(n973), .B(A[2]), .Z(n945) );
  XOR2_X2 U759 ( .A(n975), .B(A[4]), .Z(n946) );
  XOR2_X2 U760 ( .A(n977), .B(A[6]), .Z(n947) );
  XOR2_X2 U761 ( .A(A[13]), .B(A[14]), .Z(n948) );
  XOR2_X2 U762 ( .A(n983), .B(A[12]), .Z(n949) );
  XOR2_X2 U763 ( .A(n979), .B(A[8]), .Z(n950) );
  XOR2_X2 U764 ( .A(n981), .B(A[10]), .Z(n951) );
  OR2_X4 U765 ( .A1(n658), .A2(C[0]), .ZN(n952) );
  AND2_X4 U766 ( .A1(n952), .A2(n194), .ZN(MAC[0]) );
  XNOR2_X2 U767 ( .A(n51), .B(n77), .ZN(n954) );
  INV_X4 U768 ( .A(n954), .ZN(MAC[31]) );
  XNOR2_X1 U769 ( .A(A[15]), .B(B[3]), .ZN(n671) );
  XNOR2_X1 U770 ( .A(n977), .B(B[3]), .ZN(n756) );
  XNOR2_X1 U771 ( .A(n973), .B(B[3]), .ZN(n790) );
  XNOR2_X1 U772 ( .A(n975), .B(B[3]), .ZN(n773) );
  XNOR2_X1 U773 ( .A(A[13]), .B(B[3]), .ZN(n688) );
  XNOR2_X1 U774 ( .A(n979), .B(B[3]), .ZN(n739) );
  XNOR2_X1 U775 ( .A(n983), .B(B[3]), .ZN(n705) );
  XNOR2_X1 U776 ( .A(n981), .B(B[3]), .ZN(n722) );
  AOI21_X2 U777 ( .B1(n115), .B2(n956), .A(n112), .ZN(n110) );
  AOI21_X2 U778 ( .B1(n107), .B2(n957), .A(n104), .ZN(n102) );
  AOI21_X2 U779 ( .B1(n99), .B2(n958), .A(n96), .ZN(n94) );
  AOI21_X2 U780 ( .B1(n91), .B2(n959), .A(n88), .ZN(n86) );
  NAND2_X2 U781 ( .A1(n816), .A2(n966), .ZN(n18) );
  NAND2_X2 U782 ( .A1(n812), .A2(n970), .ZN(n42) );
  INV_X4 U783 ( .A(n947), .ZN(n967) );
  INV_X4 U784 ( .A(n948), .ZN(n971) );
  INV_X4 U785 ( .A(n974), .ZN(n975) );
  INV_X4 U786 ( .A(n982), .ZN(n983) );
  INV_X2 U787 ( .A(n145), .ZN(n144) );
  NOR2_X1 U788 ( .A1(n121), .A2(n124), .ZN(n119) );
  INV_X1 U789 ( .A(n148), .ZN(n209) );
  INV_X2 U790 ( .A(n143), .ZN(n141) );
  NOR2_X1 U791 ( .A1(n420), .A2(n431), .ZN(n142) );
  NAND2_X1 U792 ( .A1(n432), .A2(n441), .ZN(n149) );
  OAI22_X1 U793 ( .A1(n778), .A2(n6), .B1(n778), .B2(n834), .ZN(n512) );
  OAI22_X1 U794 ( .A1(n42), .A2(n682), .B1(n970), .B2(n681), .ZN(n546) );
  OAI22_X1 U795 ( .A1(n48), .A2(n665), .B1(n971), .B2(n664), .ZN(n529) );
  OAI21_X1 U796 ( .B1(n126), .B2(n124), .A(n125), .ZN(n123) );
  NAND2_X1 U797 ( .A1(n204), .A2(n122), .ZN(n61) );
  OAI22_X1 U798 ( .A1(n676), .A2(n42), .B1(n676), .B2(n970), .ZN(n494) );
  AOI21_X1 U799 ( .B1(n144), .B2(n135), .A(n136), .ZN(n134) );
  NAND2_X1 U800 ( .A1(n955), .A2(n133), .ZN(n63) );
  NAND2_X1 U801 ( .A1(n208), .A2(n143), .ZN(n65) );
  OAI22_X1 U802 ( .A1(n6), .A2(n791), .B1(n790), .B2(n834), .ZN(n655) );
  OAI21_X2 U803 ( .B1(n121), .B2(n125), .A(n122), .ZN(n120) );
  AOI21_X2 U804 ( .B1(n146), .B2(n154), .A(n147), .ZN(n145) );
  NOR2_X2 U805 ( .A1(n148), .A2(n151), .ZN(n146) );
  OAI21_X2 U806 ( .B1(n148), .B2(n152), .A(n149), .ZN(n147) );
  OAI21_X2 U807 ( .B1(n145), .B2(n128), .A(n129), .ZN(n127) );
  AOI21_X2 U808 ( .B1(n955), .B2(n136), .A(n131), .ZN(n129) );
  OAI21_X2 U809 ( .B1(n118), .B2(n116), .A(n117), .ZN(n115) );
  OAI21_X2 U810 ( .B1(n110), .B2(n108), .A(n109), .ZN(n107) );
  OAI21_X2 U811 ( .B1(n102), .B2(n100), .A(n101), .ZN(n99) );
  OAI21_X2 U812 ( .B1(n94), .B2(n92), .A(n93), .ZN(n91) );
  OAI21_X2 U813 ( .B1(n137), .B2(n143), .A(n138), .ZN(n136) );
  OAI21_X2 U814 ( .B1(n157), .B2(n155), .A(n156), .ZN(n154) );
  NOR2_X2 U815 ( .A1(n137), .A2(n142), .ZN(n135) );
  AOI21_X2 U816 ( .B1(n162), .B2(n963), .A(n159), .ZN(n157) );
  AOI21_X2 U817 ( .B1(n960), .B2(n180), .A(n177), .ZN(n175) );
  OAI21_X2 U818 ( .B1(n163), .B2(n175), .A(n164), .ZN(n162) );
  AOI21_X2 U819 ( .B1(n961), .B2(n171), .A(n166), .ZN(n164) );
  NOR2_X2 U820 ( .A1(n408), .A2(n419), .ZN(n137) );
  NOR2_X2 U821 ( .A1(n364), .A2(n379), .ZN(n121) );
  NOR2_X2 U822 ( .A1(n432), .A2(n441), .ZN(n148) );
  NOR2_X2 U823 ( .A1(n380), .A2(n393), .ZN(n124) );
  NOR2_X2 U824 ( .A1(n442), .A2(n451), .ZN(n151) );
  NOR2_X2 U825 ( .A1(n348), .A2(n363), .ZN(n116) );
  NOR2_X2 U826 ( .A1(n318), .A2(n331), .ZN(n108) );
  NOR2_X2 U827 ( .A1(n452), .A2(n459), .ZN(n155) );
  OR2_X1 U828 ( .A1(n394), .A2(n407), .ZN(n955) );
  OR2_X1 U829 ( .A1(n332), .A2(n347), .ZN(n956) );
  OR2_X1 U830 ( .A1(n304), .A2(n317), .ZN(n957) );
  NOR2_X2 U831 ( .A1(n292), .A2(n303), .ZN(n100) );
  NOR2_X2 U832 ( .A1(n270), .A2(n279), .ZN(n92) );
  OR2_X1 U833 ( .A1(n280), .A2(n291), .ZN(n958) );
  OR2_X1 U834 ( .A1(n260), .A2(n269), .ZN(n959) );
  NOR2_X2 U835 ( .A1(n252), .A2(n259), .ZN(n84) );
  OAI21_X2 U836 ( .B1(n181), .B2(n183), .A(n182), .ZN(n180) );
  OAI21_X2 U837 ( .B1(n86), .B2(n84), .A(n85), .ZN(n83) );
  OR2_X1 U838 ( .A1(n480), .A2(n483), .ZN(n960) );
  OR2_X1 U839 ( .A1(n468), .A2(n473), .ZN(n961) );
  OR2_X1 U840 ( .A1(n474), .A2(n479), .ZN(n962) );
  OR2_X1 U841 ( .A1(n460), .A2(n467), .ZN(n963) );
  AOI21_X2 U842 ( .B1(n964), .B2(n192), .A(n189), .ZN(n187) );
  OAI21_X2 U843 ( .B1(n187), .B2(n185), .A(n186), .ZN(n184) );
  INV_X4 U844 ( .A(n512), .ZN(n642) );
  INV_X4 U845 ( .A(n509), .ZN(n625) );
  NOR2_X2 U846 ( .A1(n484), .A2(n486), .ZN(n181) );
  INV_X4 U847 ( .A(n506), .ZN(n608) );
  NOR2_X2 U848 ( .A1(n488), .A2(n489), .ZN(n185) );
  OR2_X1 U849 ( .A1(n490), .A2(n522), .ZN(n964) );
  INV_X4 U850 ( .A(n503), .ZN(n591) );
  INV_X4 U851 ( .A(n500), .ZN(n574) );
  INV_X4 U852 ( .A(n497), .ZN(n557) );
  INV_X4 U853 ( .A(n494), .ZN(n540) );
  AOI21_X2 U854 ( .B1(n144), .B2(n208), .A(n141), .ZN(n139) );
  AOI21_X2 U855 ( .B1(n174), .B2(n962), .A(n171), .ZN(n169) );
  OAI21_X2 U856 ( .B1(n153), .B2(n151), .A(n152), .ZN(n150) );
  XNOR2_X2 U857 ( .A(C[31]), .B(n221), .ZN(n51) );
  NAND2_X2 U858 ( .A1(n815), .A2(n967), .ZN(n24) );
  NAND2_X2 U859 ( .A1(n814), .A2(n968), .ZN(n30) );
  NAND2_X2 U860 ( .A1(n813), .A2(n969), .ZN(n36) );
  NAND2_X2 U861 ( .A1(n811), .A2(n971), .ZN(n48) );
  NAND2_X2 U862 ( .A1(n817), .A2(n965), .ZN(n12) );
  NAND2_X2 U863 ( .A1(n818), .A2(n834), .ZN(n6) );
  INV_X4 U864 ( .A(A[0]), .ZN(n834) );
  INV_X4 U865 ( .A(A[15]), .ZN(n985) );
  INV_X4 U866 ( .A(n980), .ZN(n981) );
  INV_X4 U867 ( .A(A[9]), .ZN(n980) );
  INV_X4 U868 ( .A(n978), .ZN(n979) );
  INV_X4 U869 ( .A(A[7]), .ZN(n978) );
  INV_X4 U870 ( .A(n972), .ZN(n973) );
  INV_X4 U871 ( .A(A[1]), .ZN(n972) );
  INV_X4 U872 ( .A(n976), .ZN(n977) );
  INV_X4 U873 ( .A(A[5]), .ZN(n976) );
  INV_X4 U874 ( .A(A[11]), .ZN(n982) );
  INV_X4 U875 ( .A(A[3]), .ZN(n974) );
  INV_X4 U876 ( .A(n951), .ZN(n969) );
  INV_X4 U877 ( .A(n945), .ZN(n965) );
  INV_X4 U878 ( .A(n950), .ZN(n968) );
  INV_X4 U879 ( .A(n949), .ZN(n970) );
  INV_X4 U880 ( .A(n946), .ZN(n966) );
  INV_X4 U881 ( .A(n491), .ZN(n523) );
  INV_X4 U882 ( .A(n98), .ZN(n96) );
  INV_X4 U883 ( .A(n90), .ZN(n88) );
  OAI22_X2 U884 ( .A1(n761), .A2(n12), .B1(n761), .B2(n965), .ZN(n509) );
  OAI22_X2 U885 ( .A1(n744), .A2(n18), .B1(n744), .B2(n966), .ZN(n506) );
  OAI22_X2 U886 ( .A1(n727), .A2(n24), .B1(n727), .B2(n967), .ZN(n503) );
  OAI22_X2 U887 ( .A1(n710), .A2(n30), .B1(n710), .B2(n968), .ZN(n500) );
  OAI22_X2 U888 ( .A1(n693), .A2(n36), .B1(n693), .B2(n969), .ZN(n497) );
  OAI22_X2 U889 ( .A1(n659), .A2(n48), .B1(n659), .B2(n971), .ZN(n491) );
  INV_X4 U890 ( .A(C[17]), .ZN(n346) );
  INV_X4 U891 ( .A(C[19]), .ZN(n316) );
  INV_X4 U892 ( .A(C[21]), .ZN(n290) );
  INV_X4 U893 ( .A(C[23]), .ZN(n268) );
  INV_X4 U894 ( .A(C[25]), .ZN(n250) );
  INV_X4 U895 ( .A(C[27]), .ZN(n236) );
  INV_X4 U896 ( .A(C[29]), .ZN(n226) );
  INV_X4 U897 ( .A(n185), .ZN(n217) );
  INV_X4 U898 ( .A(n181), .ZN(n216) );
  INV_X4 U899 ( .A(n155), .ZN(n211) );
  INV_X4 U900 ( .A(n151), .ZN(n210) );
  INV_X4 U901 ( .A(n137), .ZN(n207) );
  INV_X4 U902 ( .A(n124), .ZN(n205) );
  INV_X4 U903 ( .A(n121), .ZN(n204) );
  INV_X4 U904 ( .A(n116), .ZN(n203) );
  INV_X4 U905 ( .A(n108), .ZN(n201) );
  INV_X4 U906 ( .A(n100), .ZN(n199) );
  INV_X4 U907 ( .A(n92), .ZN(n197) );
  INV_X4 U908 ( .A(n84), .ZN(n195) );
  INV_X4 U909 ( .A(n194), .ZN(n192) );
  INV_X4 U910 ( .A(n191), .ZN(n189) );
  INV_X4 U911 ( .A(n184), .ZN(n183) );
  INV_X4 U912 ( .A(n179), .ZN(n177) );
  INV_X4 U913 ( .A(n175), .ZN(n174) );
  INV_X4 U914 ( .A(n173), .ZN(n171) );
  INV_X4 U915 ( .A(n168), .ZN(n166) );
  INV_X4 U916 ( .A(n161), .ZN(n159) );
  INV_X4 U917 ( .A(n154), .ZN(n153) );
  INV_X4 U918 ( .A(n142), .ZN(n208) );
  INV_X4 U919 ( .A(n133), .ZN(n131) );
  INV_X4 U920 ( .A(n127), .ZN(n126) );
  INV_X4 U921 ( .A(n114), .ZN(n112) );
  INV_X4 U922 ( .A(n106), .ZN(n104) );
endmodule


module macopertion_1 ( in_a_mac, in_b_mac, bitselect1, clk, min );
  input [15:0] in_a_mac;
  input [15:0] in_b_mac;
  input [3:0] bitselect1;
  output [15:0] min;
  input clk;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18,
         N19, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49,
         N50, N51, n33, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196;
  wire   [31:0] in_c_mac;
  wire   [31:0] out_mac;
  assign min[15] = 1'b0;

  macopertion_1_DW02_mac_1 U1 ( .A(in_a_mac), .B({in_b_mac[15:1], n179}), .C(
        in_c_mac), .TC(1'b1), .MAC(out_mac) );
  SDFF_X1 in_c_mac_reg_16_ ( .D(out_mac[16]), .SI(1'b0), .SE(n33), .CK(clk), 
        .Q(in_c_mac[16]) );
  SDFF_X1 in_c_mac_reg_17_ ( .D(out_mac[17]), .SI(1'b0), .SE(n33), .CK(clk), 
        .Q(in_c_mac[17]) );
  SDFF_X1 in_c_mac_reg_18_ ( .D(out_mac[18]), .SI(1'b0), .SE(n33), .CK(clk), 
        .Q(in_c_mac[18]) );
  SDFF_X1 in_c_mac_reg_19_ ( .D(out_mac[19]), .SI(1'b0), .SE(n33), .CK(clk), 
        .Q(in_c_mac[19]) );
  SDFF_X1 in_c_mac_reg_20_ ( .D(out_mac[20]), .SI(1'b0), .SE(n33), .CK(clk), 
        .Q(in_c_mac[20]) );
  SDFF_X1 in_c_mac_reg_21_ ( .D(out_mac[21]), .SI(1'b0), .SE(n33), .CK(clk), 
        .Q(in_c_mac[21]) );
  SDFF_X1 in_c_mac_reg_22_ ( .D(out_mac[22]), .SI(1'b0), .SE(n33), .CK(clk), 
        .Q(in_c_mac[22]) );
  SDFF_X1 in_c_mac_reg_23_ ( .D(out_mac[23]), .SI(1'b0), .SE(n33), .CK(clk), 
        .Q(in_c_mac[23]) );
  SDFF_X1 in_c_mac_reg_24_ ( .D(out_mac[24]), .SI(1'b0), .SE(n33), .CK(clk), 
        .Q(in_c_mac[24]) );
  SDFF_X1 in_c_mac_reg_25_ ( .D(out_mac[25]), .SI(1'b0), .SE(n33), .CK(clk), 
        .Q(in_c_mac[25]) );
  SDFF_X1 in_c_mac_reg_26_ ( .D(out_mac[26]), .SI(1'b0), .SE(n33), .CK(clk), 
        .Q(in_c_mac[26]) );
  SDFF_X1 in_c_mac_reg_27_ ( .D(out_mac[27]), .SI(1'b0), .SE(n33), .CK(clk), 
        .Q(in_c_mac[27]) );
  SDFF_X1 in_c_mac_reg_28_ ( .D(out_mac[28]), .SI(1'b0), .SE(n33), .CK(clk), 
        .Q(in_c_mac[28]) );
  SDFF_X1 in_c_mac_reg_29_ ( .D(out_mac[29]), .SI(1'b0), .SE(n33), .CK(clk), 
        .Q(in_c_mac[29]) );
  SDFF_X1 in_c_mac_reg_30_ ( .D(out_mac[30]), .SI(1'b0), .SE(n33), .CK(clk), 
        .Q(in_c_mac[30]) );
  DFF_X1 min_reg_9_ ( .D(N46), .CK(clk), .Q(min[9]) );
  DFF_X1 min_reg_8_ ( .D(N45), .CK(clk), .Q(min[8]) );
  DFF_X1 min_reg_7_ ( .D(N44), .CK(clk), .Q(min[7]) );
  DFF_X1 min_reg_6_ ( .D(N43), .CK(clk), .Q(min[6]) );
  DFF_X1 min_reg_5_ ( .D(N42), .CK(clk), .Q(min[5]) );
  DFF_X1 min_reg_4_ ( .D(N41), .CK(clk), .Q(min[4]) );
  DFF_X1 min_reg_3_ ( .D(N40), .CK(clk), .Q(min[3]) );
  DFF_X1 min_reg_2_ ( .D(N39), .CK(clk), .Q(min[2]) );
  DFF_X1 min_reg_1_ ( .D(N38), .CK(clk), .Q(min[1]) );
  DFF_X1 min_reg_0_ ( .D(N37), .CK(clk), .Q(min[0]) );
  SDFF_X2 in_c_mac_reg_31_ ( .D(out_mac[31]), .SI(1'b0), .SE(n33), .CK(clk), 
        .Q(in_c_mac[31]) );
  DFF_X2 in_c_mac_reg_0_ ( .D(N4), .CK(clk), .Q(in_c_mac[0]) );
  DFF_X2 in_c_mac_reg_1_ ( .D(N5), .CK(clk), .Q(in_c_mac[1]) );
  DFF_X2 in_c_mac_reg_2_ ( .D(N6), .CK(clk), .Q(in_c_mac[2]) );
  DFF_X2 in_c_mac_reg_3_ ( .D(N7), .CK(clk), .Q(in_c_mac[3]) );
  DFF_X2 in_c_mac_reg_4_ ( .D(N8), .CK(clk), .Q(in_c_mac[4]) );
  DFF_X2 in_c_mac_reg_5_ ( .D(N9), .CK(clk), .Q(in_c_mac[5]) );
  DFF_X2 in_c_mac_reg_6_ ( .D(N10), .CK(clk), .Q(in_c_mac[6]) );
  DFF_X2 in_c_mac_reg_7_ ( .D(N11), .CK(clk), .Q(in_c_mac[7]) );
  DFF_X2 in_c_mac_reg_8_ ( .D(N12), .CK(clk), .Q(in_c_mac[8]) );
  DFF_X2 in_c_mac_reg_10_ ( .D(N14), .CK(clk), .Q(in_c_mac[10]) );
  DFF_X2 in_c_mac_reg_9_ ( .D(N13), .CK(clk), .Q(in_c_mac[9]) );
  DFF_X2 in_c_mac_reg_11_ ( .D(N15), .CK(clk), .Q(in_c_mac[11]) );
  DFF_X2 in_c_mac_reg_12_ ( .D(N16), .CK(clk), .Q(in_c_mac[12]) );
  DFF_X2 in_c_mac_reg_13_ ( .D(N17), .CK(clk), .Q(in_c_mac[13]) );
  DFF_X2 in_c_mac_reg_14_ ( .D(N18), .CK(clk), .Q(in_c_mac[14]) );
  DFF_X2 in_c_mac_reg_15_ ( .D(N19), .CK(clk), .Q(in_c_mac[15]) );
  DFF_X2 min_reg_14_ ( .D(N51), .CK(clk), .Q(min[14]) );
  DFF_X2 min_reg_13_ ( .D(N50), .CK(clk), .Q(min[13]) );
  DFF_X2 min_reg_12_ ( .D(N49), .CK(clk), .Q(min[12]) );
  DFF_X2 min_reg_11_ ( .D(N48), .CK(clk), .Q(min[11]) );
  DFF_X2 min_reg_10_ ( .D(N47), .CK(clk), .Q(min[10]) );
  INV_X4 U23 ( .A(n180), .ZN(n179) );
  INV_X1 U24 ( .A(in_b_mac[0]), .ZN(n180) );
  INV_X4 U25 ( .A(n181), .ZN(n33) );
  OR4_X4 U26 ( .A1(bitselect1[1]), .A2(bitselect1[0]), .A3(bitselect1[3]), 
        .A4(bitselect1[2]), .ZN(n181) );
  AND2_X1 U27 ( .A1(out_mac[15]), .A2(n181), .ZN(N19) );
  AND2_X1 U28 ( .A1(out_mac[14]), .A2(n181), .ZN(N18) );
  AND2_X1 U29 ( .A1(out_mac[13]), .A2(n181), .ZN(N17) );
  AND2_X1 U30 ( .A1(out_mac[12]), .A2(n181), .ZN(N16) );
  AND2_X1 U31 ( .A1(out_mac[11]), .A2(n181), .ZN(N15) );
  AND2_X1 U32 ( .A1(out_mac[10]), .A2(n181), .ZN(N14) );
  AND2_X1 U33 ( .A1(out_mac[9]), .A2(n181), .ZN(N13) );
  AND2_X1 U34 ( .A1(out_mac[8]), .A2(n181), .ZN(N12) );
  AND2_X1 U35 ( .A1(out_mac[7]), .A2(n181), .ZN(N11) );
  AND2_X1 U36 ( .A1(out_mac[6]), .A2(n181), .ZN(N10) );
  AND2_X1 U37 ( .A1(out_mac[5]), .A2(n181), .ZN(N9) );
  AND2_X1 U38 ( .A1(out_mac[4]), .A2(n181), .ZN(N8) );
  AND2_X1 U39 ( .A1(out_mac[3]), .A2(n181), .ZN(N7) );
  AND2_X1 U40 ( .A1(out_mac[2]), .A2(n181), .ZN(N6) );
  AND2_X1 U41 ( .A1(out_mac[1]), .A2(n181), .ZN(N5) );
  AND2_X1 U42 ( .A1(out_mac[0]), .A2(n181), .ZN(N4) );
  INV_X4 U43 ( .A(out_mac[16]), .ZN(n182) );
  NOR2_X2 U44 ( .A1(out_mac[31]), .A2(n182), .ZN(N37) );
  INV_X4 U45 ( .A(out_mac[17]), .ZN(n183) );
  NOR2_X2 U46 ( .A1(out_mac[31]), .A2(n183), .ZN(N38) );
  INV_X4 U47 ( .A(out_mac[18]), .ZN(n184) );
  NOR2_X2 U48 ( .A1(out_mac[31]), .A2(n184), .ZN(N39) );
  INV_X4 U49 ( .A(out_mac[19]), .ZN(n185) );
  NOR2_X2 U50 ( .A1(out_mac[31]), .A2(n185), .ZN(N40) );
  INV_X4 U51 ( .A(out_mac[20]), .ZN(n186) );
  NOR2_X2 U52 ( .A1(out_mac[31]), .A2(n186), .ZN(N41) );
  INV_X4 U53 ( .A(out_mac[21]), .ZN(n187) );
  NOR2_X2 U54 ( .A1(out_mac[31]), .A2(n187), .ZN(N42) );
  INV_X4 U55 ( .A(out_mac[22]), .ZN(n188) );
  NOR2_X2 U56 ( .A1(out_mac[31]), .A2(n188), .ZN(N43) );
  INV_X4 U57 ( .A(out_mac[23]), .ZN(n189) );
  NOR2_X2 U58 ( .A1(out_mac[31]), .A2(n189), .ZN(N44) );
  INV_X4 U59 ( .A(out_mac[24]), .ZN(n190) );
  NOR2_X2 U60 ( .A1(out_mac[31]), .A2(n190), .ZN(N45) );
  INV_X4 U61 ( .A(out_mac[25]), .ZN(n191) );
  NOR2_X2 U62 ( .A1(out_mac[31]), .A2(n191), .ZN(N46) );
  INV_X4 U63 ( .A(out_mac[26]), .ZN(n192) );
  NOR2_X2 U64 ( .A1(out_mac[31]), .A2(n192), .ZN(N47) );
  INV_X4 U65 ( .A(out_mac[27]), .ZN(n193) );
  NOR2_X2 U66 ( .A1(out_mac[31]), .A2(n193), .ZN(N48) );
  INV_X4 U67 ( .A(out_mac[28]), .ZN(n194) );
  NOR2_X2 U68 ( .A1(out_mac[31]), .A2(n194), .ZN(N49) );
  INV_X4 U69 ( .A(out_mac[29]), .ZN(n195) );
  NOR2_X2 U70 ( .A1(out_mac[31]), .A2(n195), .ZN(N50) );
  INV_X4 U71 ( .A(out_mac[30]), .ZN(n196) );
  NOR2_X2 U72 ( .A1(out_mac[31]), .A2(n196), .ZN(N51) );
endmodule


module macopertion_3_DW02_mac_1 ( A, B, C, TC, MAC );
  input [15:0] A;
  input [15:0] B;
  input [31:0] C;
  output [31:0] MAC;
  input TC;
  wire   n6, n12, n18, n24, n30, n36, n42, n48, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n88, n90, n91, n92, n93, n94, n96, n98, n99, n100, n101, n102,
         n104, n106, n107, n108, n109, n110, n112, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n131, n133, n134, n135, n136, n137, n138, n139, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n159, n161, n162, n163, n164, n166, n168,
         n169, n171, n173, n174, n175, n177, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n189, n191, n192, n194, n195, n197, n199,
         n201, n203, n204, n205, n207, n208, n209, n210, n211, n216, n217,
         n221, n222, n223, n224, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n494, n497, n500, n503, n506, n509, n512, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n811, n812, n813, n814, n815, n816, n817, n818, n834, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981;

  FA_X1 U53 ( .A(n223), .B(n222), .CI(n78), .CO(n77), .S(MAC[30]) );
  FA_X1 U54 ( .A(n224), .B(n227), .CI(n79), .CO(n78), .S(MAC[29]) );
  FA_X1 U55 ( .A(n231), .B(n228), .CI(n80), .CO(n79), .S(MAC[28]) );
  FA_X1 U56 ( .A(n237), .B(n232), .CI(n81), .CO(n80), .S(MAC[27]) );
  FA_X1 U58 ( .A(n244), .B(n251), .CI(n83), .CO(n82), .S(MAC[25]) );
  XOR2_X2 U59 ( .A(n52), .B(n86), .Z(MAC[24]) );
  NAND2_X2 U61 ( .A1(n195), .A2(n85), .ZN(n52) );
  NAND2_X2 U64 ( .A1(n252), .A2(n259), .ZN(n85) );
  XNOR2_X2 U65 ( .A(n91), .B(n53), .ZN(MAC[23]) );
  NAND2_X2 U69 ( .A1(n959), .A2(n90), .ZN(n53) );
  NAND2_X2 U72 ( .A1(n260), .A2(n269), .ZN(n90) );
  XOR2_X2 U73 ( .A(n54), .B(n94), .Z(MAC[22]) );
  NAND2_X2 U75 ( .A1(n197), .A2(n93), .ZN(n54) );
  NAND2_X2 U78 ( .A1(n270), .A2(n279), .ZN(n93) );
  XNOR2_X2 U79 ( .A(n99), .B(n55), .ZN(MAC[21]) );
  NAND2_X2 U83 ( .A1(n958), .A2(n98), .ZN(n55) );
  NAND2_X2 U86 ( .A1(n280), .A2(n291), .ZN(n98) );
  XOR2_X2 U87 ( .A(n56), .B(n102), .Z(MAC[20]) );
  NAND2_X2 U89 ( .A1(n199), .A2(n101), .ZN(n56) );
  NAND2_X2 U92 ( .A1(n292), .A2(n303), .ZN(n101) );
  XNOR2_X2 U93 ( .A(n107), .B(n57), .ZN(MAC[19]) );
  NAND2_X2 U97 ( .A1(n957), .A2(n106), .ZN(n57) );
  NAND2_X2 U100 ( .A1(n304), .A2(n317), .ZN(n106) );
  XOR2_X2 U101 ( .A(n58), .B(n110), .Z(MAC[18]) );
  NAND2_X2 U103 ( .A1(n201), .A2(n109), .ZN(n58) );
  NAND2_X2 U106 ( .A1(n318), .A2(n331), .ZN(n109) );
  XNOR2_X2 U107 ( .A(n115), .B(n59), .ZN(MAC[17]) );
  NAND2_X2 U111 ( .A1(n956), .A2(n114), .ZN(n59) );
  NAND2_X2 U114 ( .A1(n332), .A2(n347), .ZN(n114) );
  XOR2_X2 U115 ( .A(n60), .B(n118), .Z(MAC[16]) );
  NAND2_X2 U117 ( .A1(n203), .A2(n117), .ZN(n60) );
  NAND2_X2 U120 ( .A1(n348), .A2(n363), .ZN(n117) );
  XNOR2_X2 U121 ( .A(n123), .B(n61), .ZN(MAC[15]) );
  NAND2_X2 U128 ( .A1(n364), .A2(n379), .ZN(n122) );
  XOR2_X2 U129 ( .A(n62), .B(n126), .Z(MAC[14]) );
  NAND2_X2 U131 ( .A1(n205), .A2(n125), .ZN(n62) );
  NAND2_X2 U134 ( .A1(n380), .A2(n393), .ZN(n125) );
  XOR2_X2 U135 ( .A(n63), .B(n134), .Z(MAC[13]) );
  NAND2_X2 U138 ( .A1(n955), .A2(n135), .ZN(n128) );
  NAND2_X2 U145 ( .A1(n394), .A2(n407), .ZN(n133) );
  XOR2_X2 U146 ( .A(n64), .B(n139), .Z(MAC[12]) );
  NAND2_X2 U150 ( .A1(n207), .A2(n138), .ZN(n64) );
  NAND2_X2 U153 ( .A1(n408), .A2(n419), .ZN(n138) );
  XNOR2_X2 U154 ( .A(n144), .B(n65), .ZN(MAC[11]) );
  NAND2_X2 U161 ( .A1(n420), .A2(n431), .ZN(n143) );
  XNOR2_X2 U162 ( .A(n150), .B(n66), .ZN(MAC[10]) );
  NAND2_X2 U167 ( .A1(n209), .A2(n149), .ZN(n66) );
  XOR2_X2 U171 ( .A(n67), .B(n153), .Z(MAC[9]) );
  NAND2_X2 U173 ( .A1(n210), .A2(n152), .ZN(n67) );
  NAND2_X2 U176 ( .A1(n442), .A2(n451), .ZN(n152) );
  XOR2_X2 U177 ( .A(n157), .B(n68), .Z(MAC[8]) );
  NAND2_X2 U180 ( .A1(n211), .A2(n156), .ZN(n68) );
  NAND2_X2 U183 ( .A1(n452), .A2(n459), .ZN(n156) );
  XNOR2_X2 U184 ( .A(n69), .B(n162), .ZN(MAC[7]) );
  NAND2_X2 U188 ( .A1(n963), .A2(n161), .ZN(n69) );
  NAND2_X2 U191 ( .A1(n460), .A2(n467), .ZN(n161) );
  XOR2_X2 U192 ( .A(n70), .B(n169), .Z(MAC[6]) );
  NAND2_X2 U194 ( .A1(n961), .A2(n962), .ZN(n163) );
  NAND2_X2 U198 ( .A1(n961), .A2(n168), .ZN(n70) );
  NAND2_X2 U201 ( .A1(n468), .A2(n473), .ZN(n168) );
  XNOR2_X2 U202 ( .A(n174), .B(n71), .ZN(MAC[5]) );
  NAND2_X2 U206 ( .A1(n962), .A2(n173), .ZN(n71) );
  NAND2_X2 U209 ( .A1(n474), .A2(n479), .ZN(n173) );
  XNOR2_X2 U210 ( .A(n72), .B(n180), .ZN(MAC[4]) );
  NAND2_X2 U215 ( .A1(n960), .A2(n179), .ZN(n72) );
  NAND2_X2 U218 ( .A1(n480), .A2(n483), .ZN(n179) );
  XOR2_X2 U219 ( .A(n183), .B(n73), .Z(MAC[3]) );
  NAND2_X2 U221 ( .A1(n216), .A2(n182), .ZN(n73) );
  NAND2_X2 U224 ( .A1(n484), .A2(n486), .ZN(n182) );
  XOR2_X2 U225 ( .A(n187), .B(n74), .Z(MAC[2]) );
  NAND2_X2 U228 ( .A1(n217), .A2(n186), .ZN(n74) );
  NAND2_X2 U231 ( .A1(n488), .A2(n489), .ZN(n186) );
  XNOR2_X2 U232 ( .A(n75), .B(n192), .ZN(MAC[1]) );
  NAND2_X2 U236 ( .A1(n964), .A2(n191), .ZN(n75) );
  NAND2_X2 U239 ( .A1(n490), .A2(n522), .ZN(n191) );
  NAND2_X2 U245 ( .A1(n658), .A2(C[0]), .ZN(n194) );
  FA_X1 U247 ( .A(C[29]), .B(C[30]), .CI(n523), .CO(n221), .S(n222) );
  FA_X1 U248 ( .A(n524), .B(n226), .CI(n229), .CO(n223), .S(n224) );
  FA_X1 U250 ( .A(n233), .B(n540), .CI(n230), .CO(n227), .S(n228) );
  FA_X1 U251 ( .A(C[27]), .B(C[28]), .CI(n525), .CO(n229), .S(n230) );
  FA_X1 U252 ( .A(n234), .B(n241), .CI(n239), .CO(n231), .S(n232) );
  FA_X1 U253 ( .A(n541), .B(n236), .CI(n526), .CO(n233), .S(n234) );
  FA_X1 U255 ( .A(n245), .B(n242), .CI(n240), .CO(n237), .S(n238) );
  FA_X1 U256 ( .A(n557), .B(n527), .CI(n247), .CO(n239), .S(n240) );
  FA_X1 U257 ( .A(C[25]), .B(C[26]), .CI(n542), .CO(n241), .S(n242) );
  FA_X1 U258 ( .A(n246), .B(n248), .CI(n253), .CO(n243), .S(n244) );
  FA_X1 U259 ( .A(n257), .B(n528), .CI(n255), .CO(n245), .S(n246) );
  FA_X1 U260 ( .A(n558), .B(n250), .CI(n543), .CO(n247), .S(n248) );
  FA_X1 U262 ( .A(n254), .B(n263), .CI(n261), .CO(n251), .S(n252) );
  FA_X1 U263 ( .A(n258), .B(n265), .CI(n256), .CO(n253), .S(n254) );
  FA_X1 U264 ( .A(n544), .B(n529), .CI(n574), .CO(n255), .S(n256) );
  FA_X1 U265 ( .A(C[23]), .B(C[24]), .CI(n559), .CO(n257), .S(n258) );
  FA_X1 U266 ( .A(n271), .B(n264), .CI(n262), .CO(n259), .S(n260) );
  FA_X1 U267 ( .A(n266), .B(n275), .CI(n273), .CO(n261), .S(n262) );
  FA_X1 U268 ( .A(n530), .B(n545), .CI(n277), .CO(n263), .S(n264) );
  FA_X1 U269 ( .A(n575), .B(n268), .CI(n560), .CO(n265), .S(n266) );
  FA_X1 U271 ( .A(n281), .B(n274), .CI(n272), .CO(n269), .S(n270) );
  FA_X1 U272 ( .A(n276), .B(n278), .CI(n283), .CO(n271), .S(n272) );
  FA_X1 U273 ( .A(n287), .B(n576), .CI(n285), .CO(n273), .S(n274) );
  FA_X1 U274 ( .A(n531), .B(n546), .CI(n591), .CO(n275), .S(n276) );
  FA_X1 U275 ( .A(C[21]), .B(C[22]), .CI(n561), .CO(n277), .S(n278) );
  FA_X1 U276 ( .A(n293), .B(n284), .CI(n282), .CO(n279), .S(n280) );
  FA_X1 U277 ( .A(n297), .B(n286), .CI(n295), .CO(n281), .S(n282) );
  FA_X1 U278 ( .A(n299), .B(n301), .CI(n288), .CO(n283), .S(n284) );
  FA_X1 U279 ( .A(n547), .B(n532), .CI(n562), .CO(n285), .S(n286) );
  FA_X1 U280 ( .A(n592), .B(n290), .CI(n577), .CO(n287), .S(n288) );
  FA_X1 U282 ( .A(n305), .B(n296), .CI(n294), .CO(n291), .S(n292) );
  FA_X1 U283 ( .A(n298), .B(n309), .CI(n307), .CO(n293), .S(n294) );
  FA_X1 U284 ( .A(n302), .B(n311), .CI(n300), .CO(n295), .S(n296) );
  FA_X1 U285 ( .A(n533), .B(n548), .CI(n313), .CO(n297), .S(n298) );
  FA_X1 U286 ( .A(n593), .B(n563), .CI(n608), .CO(n299), .S(n300) );
  FA_X1 U287 ( .A(C[19]), .B(C[20]), .CI(n578), .CO(n301), .S(n302) );
  FA_X1 U288 ( .A(n319), .B(n308), .CI(n306), .CO(n303), .S(n304) );
  FA_X1 U289 ( .A(n310), .B(n323), .CI(n321), .CO(n305), .S(n306) );
  FA_X1 U290 ( .A(n314), .B(n325), .CI(n312), .CO(n307), .S(n308) );
  FA_X1 U291 ( .A(n329), .B(n549), .CI(n327), .CO(n309), .S(n310) );
  FA_X1 U292 ( .A(n534), .B(n579), .CI(n564), .CO(n311), .S(n312) );
  FA_X1 U293 ( .A(n609), .B(n316), .CI(n594), .CO(n313), .S(n314) );
  FA_X1 U295 ( .A(n333), .B(n322), .CI(n320), .CO(n317), .S(n318) );
  FA_X1 U296 ( .A(n324), .B(n337), .CI(n335), .CO(n319), .S(n320) );
  FA_X1 U297 ( .A(n326), .B(n330), .CI(n328), .CO(n321), .S(n322) );
  FA_X1 U298 ( .A(n341), .B(n343), .CI(n339), .CO(n323), .S(n324) );
  FA_X1 U299 ( .A(n550), .B(n610), .CI(n595), .CO(n325), .S(n326) );
  FA_X1 U300 ( .A(n535), .B(n565), .CI(n625), .CO(n327), .S(n328) );
  FA_X1 U301 ( .A(C[17]), .B(C[18]), .CI(n580), .CO(n329), .S(n330) );
  FA_X1 U302 ( .A(n349), .B(n336), .CI(n334), .CO(n331), .S(n332) );
  FA_X1 U303 ( .A(n338), .B(n353), .CI(n351), .CO(n333), .S(n334) );
  FA_X1 U304 ( .A(n342), .B(n344), .CI(n340), .CO(n335), .S(n336) );
  FA_X1 U305 ( .A(n357), .B(n359), .CI(n355), .CO(n337), .S(n338) );
  FA_X1 U306 ( .A(n566), .B(n581), .CI(n361), .CO(n339), .S(n340) );
  FA_X1 U307 ( .A(n536), .B(n596), .CI(n551), .CO(n341), .S(n342) );
  FA_X1 U308 ( .A(n626), .B(n346), .CI(n611), .CO(n343), .S(n344) );
  FA_X1 U310 ( .A(n365), .B(n352), .CI(n350), .CO(n347), .S(n348) );
  FA_X1 U311 ( .A(n354), .B(n369), .CI(n367), .CO(n349), .S(n350) );
  FA_X1 U312 ( .A(n371), .B(n360), .CI(n356), .CO(n351), .S(n352) );
  FA_X1 U313 ( .A(n373), .B(n375), .CI(n358), .CO(n353), .S(n354) );
  FA_X1 U314 ( .A(n377), .B(n582), .CI(n362), .CO(n355), .S(n356) );
  FA_X1 U315 ( .A(n537), .B(n612), .CI(n552), .CO(n357), .S(n358) );
  FA_X1 U316 ( .A(n627), .B(n567), .CI(n642), .CO(n359), .S(n360) );
  XNOR2_X2 U317 ( .A(n597), .B(C[16]), .ZN(n362) );
  OR2_X2 U318 ( .A1(n597), .A2(C[16]), .ZN(n361) );
  FA_X1 U319 ( .A(n381), .B(n368), .CI(n366), .CO(n363), .S(n364) );
  FA_X1 U320 ( .A(n383), .B(n372), .CI(n370), .CO(n365), .S(n366) );
  FA_X1 U321 ( .A(n376), .B(n374), .CI(n385), .CO(n367), .S(n368) );
  FA_X1 U322 ( .A(n389), .B(n378), .CI(n387), .CO(n369), .S(n370) );
  FA_X1 U323 ( .A(n598), .B(n613), .CI(n391), .CO(n371), .S(n372) );
  FA_X1 U324 ( .A(n553), .B(n568), .CI(n583), .CO(n373), .S(n374) );
  FA_X1 U325 ( .A(n515), .B(n643), .CI(n628), .CO(n375), .S(n376) );
  HA_X1 U326 ( .A(C[15]), .B(n538), .CO(n377), .S(n378) );
  FA_X1 U327 ( .A(n395), .B(n384), .CI(n382), .CO(n379), .S(n380) );
  FA_X1 U328 ( .A(n397), .B(n399), .CI(n386), .CO(n381), .S(n382) );
  FA_X1 U330 ( .A(n403), .B(n405), .CI(n401), .CO(n385), .S(n386) );
  FA_X1 U331 ( .A(n584), .B(n614), .CI(n599), .CO(n387), .S(n388) );
  FA_X1 U332 ( .A(n554), .B(n629), .CI(n569), .CO(n389), .S(n390) );
  FA_X1 U333 ( .A(n539), .B(C[14]), .CI(n644), .CO(n391), .S(n392) );
  FA_X1 U334 ( .A(n398), .B(n409), .CI(n396), .CO(n393), .S(n394) );
  FA_X1 U335 ( .A(n411), .B(n404), .CI(n400), .CO(n395), .S(n396) );
  FA_X1 U336 ( .A(n413), .B(n415), .CI(n402), .CO(n397), .S(n398) );
  FA_X1 U337 ( .A(n417), .B(n615), .CI(n406), .CO(n399), .S(n400) );
  FA_X1 U338 ( .A(n630), .B(n585), .CI(n600), .CO(n401), .S(n402) );
  FA_X1 U339 ( .A(n516), .B(n645), .CI(n570), .CO(n403), .S(n404) );
  HA_X1 U340 ( .A(C[13]), .B(n555), .CO(n405), .S(n406) );
  FA_X1 U341 ( .A(n421), .B(n412), .CI(n410), .CO(n407), .S(n408) );
  FA_X1 U342 ( .A(n414), .B(n416), .CI(n423), .CO(n409), .S(n410) );
  FA_X1 U343 ( .A(n425), .B(n427), .CI(n418), .CO(n411), .S(n412) );
  FA_X1 U344 ( .A(n601), .B(n616), .CI(n429), .CO(n413), .S(n414) );
  FA_X1 U345 ( .A(n571), .B(n631), .CI(n586), .CO(n415), .S(n416) );
  FA_X1 U346 ( .A(n556), .B(C[12]), .CI(n646), .CO(n417), .S(n418) );
  FA_X1 U347 ( .A(n433), .B(n424), .CI(n422), .CO(n419), .S(n420) );
  FA_X1 U348 ( .A(n428), .B(n426), .CI(n435), .CO(n421), .S(n422) );
  FA_X1 U349 ( .A(n430), .B(n439), .CI(n437), .CO(n423), .S(n424) );
  FA_X1 U350 ( .A(n587), .B(n617), .CI(n602), .CO(n425), .S(n426) );
  FA_X1 U351 ( .A(n517), .B(n647), .CI(n632), .CO(n427), .S(n428) );
  HA_X1 U352 ( .A(C[11]), .B(n572), .CO(n429), .S(n430) );
  FA_X1 U353 ( .A(n443), .B(n436), .CI(n434), .CO(n431), .S(n432) );
  FA_X1 U354 ( .A(n438), .B(n440), .CI(n445), .CO(n433), .S(n434) );
  FA_X1 U355 ( .A(n449), .B(n618), .CI(n447), .CO(n435), .S(n436) );
  FA_X1 U356 ( .A(n588), .B(n633), .CI(n603), .CO(n437), .S(n438) );
  FA_X1 U357 ( .A(n573), .B(C[10]), .CI(n648), .CO(n439), .S(n440) );
  FA_X1 U358 ( .A(n453), .B(n446), .CI(n444), .CO(n441), .S(n442) );
  FA_X1 U359 ( .A(n455), .B(n450), .CI(n448), .CO(n443), .S(n444) );
  FA_X1 U360 ( .A(n604), .B(n619), .CI(n457), .CO(n445), .S(n446) );
  FA_X1 U361 ( .A(n518), .B(n649), .CI(n634), .CO(n447), .S(n448) );
  HA_X1 U362 ( .A(C[9]), .B(n589), .CO(n449), .S(n450) );
  FA_X1 U363 ( .A(n461), .B(n456), .CI(n454), .CO(n451), .S(n452) );
  FA_X1 U364 ( .A(n463), .B(n465), .CI(n458), .CO(n453), .S(n454) );
  FA_X1 U365 ( .A(n605), .B(n635), .CI(n620), .CO(n455), .S(n456) );
  FA_X1 U366 ( .A(n590), .B(C[8]), .CI(n650), .CO(n457), .S(n458) );
  FA_X1 U367 ( .A(n464), .B(n469), .CI(n462), .CO(n459), .S(n460) );
  FA_X1 U368 ( .A(n471), .B(n636), .CI(n466), .CO(n461), .S(n462) );
  FA_X1 U369 ( .A(n519), .B(n651), .CI(n621), .CO(n463), .S(n464) );
  HA_X1 U370 ( .A(C[7]), .B(n606), .CO(n465), .S(n466) );
  FA_X1 U371 ( .A(n472), .B(n475), .CI(n470), .CO(n467), .S(n468) );
  FA_X1 U372 ( .A(n622), .B(n637), .CI(n477), .CO(n469), .S(n470) );
  FA_X1 U373 ( .A(n607), .B(C[6]), .CI(n652), .CO(n471), .S(n472) );
  FA_X1 U374 ( .A(n478), .B(n481), .CI(n476), .CO(n473), .S(n474) );
  FA_X1 U375 ( .A(n520), .B(n653), .CI(n638), .CO(n475), .S(n476) );
  HA_X1 U376 ( .A(C[5]), .B(n623), .CO(n477), .S(n478) );
  FA_X1 U377 ( .A(n485), .B(n639), .CI(n482), .CO(n479), .S(n480) );
  FA_X1 U378 ( .A(n624), .B(C[4]), .CI(n654), .CO(n481), .S(n482) );
  FA_X1 U379 ( .A(n521), .B(n640), .CI(n487), .CO(n483), .S(n484) );
  HA_X1 U380 ( .A(C[3]), .B(n655), .CO(n485), .S(n486) );
  FA_X1 U381 ( .A(n641), .B(C[2]), .CI(n656), .CO(n487), .S(n488) );
  HA_X1 U382 ( .A(C[1]), .B(n657), .CO(n489), .S(n490) );
  OAI22_X2 U383 ( .A1(n48), .A2(n981), .B1(n675), .B2(n971), .ZN(n515) );
  OAI22_X2 U386 ( .A1(n48), .A2(n660), .B1(n971), .B2(n659), .ZN(n524) );
  OAI22_X2 U387 ( .A1(n48), .A2(n661), .B1(n971), .B2(n660), .ZN(n525) );
  OAI22_X2 U388 ( .A1(n48), .A2(n662), .B1(n971), .B2(n661), .ZN(n526) );
  OAI22_X2 U389 ( .A1(n48), .A2(n663), .B1(n971), .B2(n662), .ZN(n527) );
  OAI22_X2 U390 ( .A1(n48), .A2(n664), .B1(n971), .B2(n663), .ZN(n528) );
  OAI22_X2 U392 ( .A1(n48), .A2(n666), .B1(n971), .B2(n665), .ZN(n530) );
  OAI22_X2 U393 ( .A1(n48), .A2(n667), .B1(n971), .B2(n666), .ZN(n531) );
  OAI22_X2 U394 ( .A1(n48), .A2(n668), .B1(n971), .B2(n667), .ZN(n532) );
  OAI22_X2 U395 ( .A1(n48), .A2(n669), .B1(n971), .B2(n668), .ZN(n533) );
  OAI22_X2 U396 ( .A1(n48), .A2(n670), .B1(n971), .B2(n669), .ZN(n534) );
  OAI22_X2 U397 ( .A1(n48), .A2(n671), .B1(n971), .B2(n670), .ZN(n535) );
  OAI22_X2 U398 ( .A1(n48), .A2(n672), .B1(n971), .B2(n671), .ZN(n536) );
  OAI22_X2 U399 ( .A1(n48), .A2(n673), .B1(n971), .B2(n672), .ZN(n537) );
  OAI22_X2 U400 ( .A1(n48), .A2(n674), .B1(n971), .B2(n673), .ZN(n538) );
  AND2_X2 U401 ( .A1(B[0]), .A2(n946), .ZN(n539) );
  XNOR2_X2 U403 ( .A(A[15]), .B(B[15]), .ZN(n659) );
  XNOR2_X2 U404 ( .A(A[15]), .B(B[14]), .ZN(n660) );
  XNOR2_X2 U405 ( .A(A[15]), .B(B[13]), .ZN(n661) );
  XNOR2_X2 U406 ( .A(A[15]), .B(B[12]), .ZN(n662) );
  XNOR2_X2 U407 ( .A(A[15]), .B(B[11]), .ZN(n663) );
  XNOR2_X2 U408 ( .A(A[15]), .B(B[10]), .ZN(n664) );
  XNOR2_X2 U409 ( .A(A[15]), .B(B[9]), .ZN(n665) );
  XNOR2_X2 U410 ( .A(A[15]), .B(B[8]), .ZN(n666) );
  XNOR2_X2 U411 ( .A(A[15]), .B(B[7]), .ZN(n667) );
  XNOR2_X2 U412 ( .A(A[15]), .B(B[6]), .ZN(n668) );
  XNOR2_X2 U413 ( .A(A[15]), .B(B[5]), .ZN(n669) );
  XNOR2_X2 U414 ( .A(A[15]), .B(B[4]), .ZN(n670) );
  XNOR2_X2 U416 ( .A(A[15]), .B(B[2]), .ZN(n672) );
  XNOR2_X2 U417 ( .A(A[15]), .B(B[1]), .ZN(n673) );
  XNOR2_X2 U418 ( .A(B[0]), .B(A[15]), .ZN(n674) );
  OR2_X2 U419 ( .A1(B[0]), .A2(n981), .ZN(n675) );
  OAI22_X2 U421 ( .A1(n42), .A2(n980), .B1(n692), .B2(n970), .ZN(n516) );
  OAI22_X2 U424 ( .A1(n42), .A2(n677), .B1(n970), .B2(n676), .ZN(n541) );
  OAI22_X2 U425 ( .A1(n42), .A2(n678), .B1(n970), .B2(n677), .ZN(n542) );
  OAI22_X2 U426 ( .A1(n42), .A2(n679), .B1(n970), .B2(n678), .ZN(n543) );
  OAI22_X2 U427 ( .A1(n42), .A2(n680), .B1(n970), .B2(n679), .ZN(n544) );
  OAI22_X2 U428 ( .A1(n42), .A2(n681), .B1(n970), .B2(n680), .ZN(n545) );
  OAI22_X2 U430 ( .A1(n42), .A2(n683), .B1(n970), .B2(n682), .ZN(n547) );
  OAI22_X2 U431 ( .A1(n42), .A2(n684), .B1(n970), .B2(n683), .ZN(n548) );
  OAI22_X2 U432 ( .A1(n42), .A2(n685), .B1(n970), .B2(n684), .ZN(n549) );
  OAI22_X2 U433 ( .A1(n42), .A2(n686), .B1(n970), .B2(n685), .ZN(n550) );
  OAI22_X2 U434 ( .A1(n42), .A2(n687), .B1(n970), .B2(n686), .ZN(n551) );
  OAI22_X2 U435 ( .A1(n42), .A2(n688), .B1(n970), .B2(n687), .ZN(n552) );
  OAI22_X2 U436 ( .A1(n42), .A2(n689), .B1(n970), .B2(n688), .ZN(n553) );
  OAI22_X2 U437 ( .A1(n42), .A2(n690), .B1(n970), .B2(n689), .ZN(n554) );
  OAI22_X2 U438 ( .A1(n42), .A2(n691), .B1(n970), .B2(n690), .ZN(n555) );
  AND2_X2 U439 ( .A1(B[0]), .A2(n947), .ZN(n556) );
  XNOR2_X2 U441 ( .A(A[13]), .B(B[15]), .ZN(n676) );
  XNOR2_X2 U442 ( .A(A[13]), .B(B[14]), .ZN(n677) );
  XNOR2_X2 U443 ( .A(A[13]), .B(B[13]), .ZN(n678) );
  XNOR2_X2 U444 ( .A(A[13]), .B(B[12]), .ZN(n679) );
  XNOR2_X2 U445 ( .A(A[13]), .B(B[11]), .ZN(n680) );
  XNOR2_X2 U446 ( .A(A[13]), .B(B[10]), .ZN(n681) );
  XNOR2_X2 U447 ( .A(A[13]), .B(B[9]), .ZN(n682) );
  XNOR2_X2 U448 ( .A(A[13]), .B(B[8]), .ZN(n683) );
  XNOR2_X2 U449 ( .A(A[13]), .B(B[7]), .ZN(n684) );
  XNOR2_X2 U450 ( .A(A[13]), .B(B[6]), .ZN(n685) );
  XNOR2_X2 U451 ( .A(A[13]), .B(B[5]), .ZN(n686) );
  XNOR2_X2 U452 ( .A(A[13]), .B(B[4]), .ZN(n687) );
  XNOR2_X2 U454 ( .A(A[13]), .B(B[2]), .ZN(n689) );
  XNOR2_X2 U455 ( .A(A[13]), .B(B[1]), .ZN(n690) );
  XNOR2_X2 U456 ( .A(B[0]), .B(A[13]), .ZN(n691) );
  OR2_X2 U457 ( .A1(B[0]), .A2(n980), .ZN(n692) );
  OAI22_X2 U459 ( .A1(n36), .A2(n978), .B1(n709), .B2(n969), .ZN(n517) );
  OAI22_X2 U462 ( .A1(n36), .A2(n694), .B1(n969), .B2(n693), .ZN(n558) );
  OAI22_X2 U463 ( .A1(n36), .A2(n695), .B1(n969), .B2(n694), .ZN(n559) );
  OAI22_X2 U464 ( .A1(n36), .A2(n696), .B1(n969), .B2(n695), .ZN(n560) );
  OAI22_X2 U465 ( .A1(n36), .A2(n697), .B1(n969), .B2(n696), .ZN(n561) );
  OAI22_X2 U466 ( .A1(n36), .A2(n698), .B1(n969), .B2(n697), .ZN(n562) );
  OAI22_X2 U467 ( .A1(n36), .A2(n699), .B1(n969), .B2(n698), .ZN(n563) );
  OAI22_X2 U468 ( .A1(n36), .A2(n700), .B1(n969), .B2(n699), .ZN(n564) );
  OAI22_X2 U469 ( .A1(n36), .A2(n701), .B1(n969), .B2(n700), .ZN(n565) );
  OAI22_X2 U470 ( .A1(n36), .A2(n702), .B1(n969), .B2(n701), .ZN(n566) );
  OAI22_X2 U471 ( .A1(n36), .A2(n703), .B1(n969), .B2(n702), .ZN(n567) );
  OAI22_X2 U472 ( .A1(n36), .A2(n704), .B1(n969), .B2(n703), .ZN(n568) );
  OAI22_X2 U473 ( .A1(n36), .A2(n705), .B1(n969), .B2(n704), .ZN(n569) );
  OAI22_X2 U474 ( .A1(n36), .A2(n706), .B1(n969), .B2(n705), .ZN(n570) );
  OAI22_X2 U475 ( .A1(n36), .A2(n707), .B1(n969), .B2(n706), .ZN(n571) );
  OAI22_X2 U476 ( .A1(n36), .A2(n708), .B1(n969), .B2(n707), .ZN(n572) );
  AND2_X2 U477 ( .A1(B[0]), .A2(n951), .ZN(n573) );
  XNOR2_X2 U479 ( .A(n979), .B(B[15]), .ZN(n693) );
  XNOR2_X2 U480 ( .A(n979), .B(B[14]), .ZN(n694) );
  XNOR2_X2 U481 ( .A(n979), .B(B[13]), .ZN(n695) );
  XNOR2_X2 U482 ( .A(n979), .B(B[12]), .ZN(n696) );
  XNOR2_X2 U483 ( .A(n979), .B(B[11]), .ZN(n697) );
  XNOR2_X2 U484 ( .A(n979), .B(B[10]), .ZN(n698) );
  XNOR2_X2 U485 ( .A(n979), .B(B[9]), .ZN(n699) );
  XNOR2_X2 U486 ( .A(n979), .B(B[8]), .ZN(n700) );
  XNOR2_X2 U487 ( .A(n979), .B(B[7]), .ZN(n701) );
  XNOR2_X2 U488 ( .A(n979), .B(B[6]), .ZN(n702) );
  XNOR2_X2 U489 ( .A(n979), .B(B[5]), .ZN(n703) );
  XNOR2_X2 U490 ( .A(n979), .B(B[4]), .ZN(n704) );
  XNOR2_X2 U492 ( .A(n979), .B(B[2]), .ZN(n706) );
  XNOR2_X2 U493 ( .A(n979), .B(B[1]), .ZN(n707) );
  XNOR2_X2 U494 ( .A(B[0]), .B(n979), .ZN(n708) );
  OR2_X2 U495 ( .A1(B[0]), .A2(n978), .ZN(n709) );
  OAI22_X2 U497 ( .A1(n30), .A2(n977), .B1(n726), .B2(n968), .ZN(n518) );
  OAI22_X2 U500 ( .A1(n30), .A2(n711), .B1(n968), .B2(n710), .ZN(n575) );
  OAI22_X2 U501 ( .A1(n30), .A2(n712), .B1(n968), .B2(n711), .ZN(n576) );
  OAI22_X2 U502 ( .A1(n30), .A2(n713), .B1(n968), .B2(n712), .ZN(n577) );
  OAI22_X2 U503 ( .A1(n30), .A2(n714), .B1(n968), .B2(n713), .ZN(n578) );
  OAI22_X2 U504 ( .A1(n30), .A2(n715), .B1(n968), .B2(n714), .ZN(n579) );
  OAI22_X2 U505 ( .A1(n30), .A2(n716), .B1(n968), .B2(n715), .ZN(n580) );
  OAI22_X2 U506 ( .A1(n30), .A2(n717), .B1(n968), .B2(n716), .ZN(n581) );
  OAI22_X2 U507 ( .A1(n30), .A2(n718), .B1(n968), .B2(n717), .ZN(n582) );
  OAI22_X2 U508 ( .A1(n30), .A2(n719), .B1(n968), .B2(n718), .ZN(n583) );
  OAI22_X2 U509 ( .A1(n30), .A2(n720), .B1(n968), .B2(n719), .ZN(n584) );
  OAI22_X2 U510 ( .A1(n30), .A2(n721), .B1(n968), .B2(n720), .ZN(n585) );
  OAI22_X2 U511 ( .A1(n30), .A2(n722), .B1(n968), .B2(n721), .ZN(n586) );
  OAI22_X2 U512 ( .A1(n30), .A2(n723), .B1(n968), .B2(n722), .ZN(n587) );
  OAI22_X2 U513 ( .A1(n30), .A2(n724), .B1(n968), .B2(n723), .ZN(n588) );
  OAI22_X2 U514 ( .A1(n30), .A2(n725), .B1(n968), .B2(n724), .ZN(n589) );
  AND2_X2 U515 ( .A1(B[0]), .A2(n950), .ZN(n590) );
  XNOR2_X2 U517 ( .A(A[9]), .B(B[15]), .ZN(n710) );
  XNOR2_X2 U518 ( .A(A[9]), .B(B[14]), .ZN(n711) );
  XNOR2_X2 U519 ( .A(A[9]), .B(B[13]), .ZN(n712) );
  XNOR2_X2 U520 ( .A(A[9]), .B(B[12]), .ZN(n713) );
  XNOR2_X2 U521 ( .A(A[9]), .B(B[11]), .ZN(n714) );
  XNOR2_X2 U522 ( .A(A[9]), .B(B[10]), .ZN(n715) );
  XNOR2_X2 U523 ( .A(A[9]), .B(B[9]), .ZN(n716) );
  XNOR2_X2 U524 ( .A(A[9]), .B(B[8]), .ZN(n717) );
  XNOR2_X2 U525 ( .A(A[9]), .B(B[7]), .ZN(n718) );
  XNOR2_X2 U526 ( .A(A[9]), .B(B[6]), .ZN(n719) );
  XNOR2_X2 U527 ( .A(A[9]), .B(B[5]), .ZN(n720) );
  XNOR2_X2 U528 ( .A(A[9]), .B(B[4]), .ZN(n721) );
  XNOR2_X2 U530 ( .A(A[9]), .B(B[2]), .ZN(n723) );
  XNOR2_X2 U531 ( .A(A[9]), .B(B[1]), .ZN(n724) );
  XNOR2_X2 U532 ( .A(B[0]), .B(A[9]), .ZN(n725) );
  OR2_X2 U533 ( .A1(B[0]), .A2(n977), .ZN(n726) );
  OAI22_X2 U535 ( .A1(n24), .A2(n976), .B1(n743), .B2(n967), .ZN(n519) );
  OAI22_X2 U538 ( .A1(n24), .A2(n728), .B1(n967), .B2(n727), .ZN(n592) );
  OAI22_X2 U539 ( .A1(n24), .A2(n729), .B1(n967), .B2(n728), .ZN(n593) );
  OAI22_X2 U540 ( .A1(n24), .A2(n730), .B1(n967), .B2(n729), .ZN(n594) );
  OAI22_X2 U541 ( .A1(n24), .A2(n731), .B1(n967), .B2(n730), .ZN(n595) );
  OAI22_X2 U542 ( .A1(n24), .A2(n732), .B1(n967), .B2(n731), .ZN(n596) );
  OAI22_X2 U543 ( .A1(n24), .A2(n733), .B1(n967), .B2(n732), .ZN(n597) );
  OAI22_X2 U544 ( .A1(n24), .A2(n734), .B1(n967), .B2(n733), .ZN(n598) );
  OAI22_X2 U545 ( .A1(n24), .A2(n735), .B1(n967), .B2(n734), .ZN(n599) );
  OAI22_X2 U546 ( .A1(n24), .A2(n736), .B1(n967), .B2(n735), .ZN(n600) );
  OAI22_X2 U547 ( .A1(n24), .A2(n737), .B1(n967), .B2(n736), .ZN(n601) );
  OAI22_X2 U548 ( .A1(n24), .A2(n738), .B1(n967), .B2(n737), .ZN(n602) );
  OAI22_X2 U549 ( .A1(n24), .A2(n739), .B1(n967), .B2(n738), .ZN(n603) );
  OAI22_X2 U550 ( .A1(n24), .A2(n740), .B1(n967), .B2(n739), .ZN(n604) );
  OAI22_X2 U551 ( .A1(n24), .A2(n741), .B1(n967), .B2(n740), .ZN(n605) );
  OAI22_X2 U552 ( .A1(n24), .A2(n742), .B1(n967), .B2(n741), .ZN(n606) );
  AND2_X2 U553 ( .A1(B[0]), .A2(n945), .ZN(n607) );
  XNOR2_X2 U555 ( .A(A[7]), .B(B[15]), .ZN(n727) );
  XNOR2_X2 U556 ( .A(A[7]), .B(B[14]), .ZN(n728) );
  XNOR2_X2 U557 ( .A(A[7]), .B(B[13]), .ZN(n729) );
  XNOR2_X2 U558 ( .A(A[7]), .B(B[12]), .ZN(n730) );
  XNOR2_X2 U559 ( .A(A[7]), .B(B[11]), .ZN(n731) );
  XNOR2_X2 U560 ( .A(A[7]), .B(B[10]), .ZN(n732) );
  XNOR2_X2 U561 ( .A(A[7]), .B(B[9]), .ZN(n733) );
  XNOR2_X2 U564 ( .A(A[7]), .B(B[6]), .ZN(n736) );
  XNOR2_X2 U566 ( .A(A[7]), .B(B[4]), .ZN(n738) );
  XNOR2_X2 U568 ( .A(A[7]), .B(B[2]), .ZN(n740) );
  XNOR2_X2 U569 ( .A(A[7]), .B(B[1]), .ZN(n741) );
  XNOR2_X2 U570 ( .A(B[0]), .B(A[7]), .ZN(n742) );
  OR2_X2 U571 ( .A1(B[0]), .A2(n976), .ZN(n743) );
  OAI22_X2 U573 ( .A1(n18), .A2(n975), .B1(n760), .B2(n966), .ZN(n520) );
  OAI22_X2 U576 ( .A1(n18), .A2(n745), .B1(n966), .B2(n744), .ZN(n609) );
  OAI22_X2 U577 ( .A1(n18), .A2(n746), .B1(n966), .B2(n745), .ZN(n610) );
  OAI22_X2 U578 ( .A1(n18), .A2(n747), .B1(n966), .B2(n746), .ZN(n611) );
  OAI22_X2 U579 ( .A1(n18), .A2(n748), .B1(n966), .B2(n747), .ZN(n612) );
  OAI22_X2 U580 ( .A1(n18), .A2(n749), .B1(n966), .B2(n748), .ZN(n613) );
  OAI22_X2 U581 ( .A1(n18), .A2(n750), .B1(n966), .B2(n749), .ZN(n614) );
  OAI22_X2 U582 ( .A1(n18), .A2(n751), .B1(n966), .B2(n750), .ZN(n615) );
  OAI22_X2 U583 ( .A1(n18), .A2(n752), .B1(n966), .B2(n751), .ZN(n616) );
  OAI22_X2 U584 ( .A1(n18), .A2(n753), .B1(n966), .B2(n752), .ZN(n617) );
  OAI22_X2 U585 ( .A1(n18), .A2(n754), .B1(n966), .B2(n753), .ZN(n618) );
  OAI22_X2 U586 ( .A1(n18), .A2(n755), .B1(n966), .B2(n754), .ZN(n619) );
  OAI22_X2 U587 ( .A1(n18), .A2(n756), .B1(n966), .B2(n755), .ZN(n620) );
  OAI22_X2 U588 ( .A1(n18), .A2(n757), .B1(n966), .B2(n756), .ZN(n621) );
  OAI22_X2 U589 ( .A1(n18), .A2(n758), .B1(n966), .B2(n757), .ZN(n622) );
  OAI22_X2 U590 ( .A1(n18), .A2(n759), .B1(n966), .B2(n758), .ZN(n623) );
  AND2_X2 U591 ( .A1(B[0]), .A2(n949), .ZN(n624) );
  XNOR2_X2 U594 ( .A(A[5]), .B(B[14]), .ZN(n745) );
  XNOR2_X2 U595 ( .A(A[5]), .B(B[13]), .ZN(n746) );
  XNOR2_X2 U596 ( .A(A[5]), .B(B[12]), .ZN(n747) );
  XNOR2_X2 U597 ( .A(A[5]), .B(B[11]), .ZN(n748) );
  XNOR2_X2 U598 ( .A(A[5]), .B(B[10]), .ZN(n749) );
  XNOR2_X2 U599 ( .A(A[5]), .B(B[9]), .ZN(n750) );
  XNOR2_X2 U600 ( .A(A[5]), .B(B[8]), .ZN(n751) );
  XNOR2_X2 U601 ( .A(A[5]), .B(B[7]), .ZN(n752) );
  XNOR2_X2 U602 ( .A(A[5]), .B(B[6]), .ZN(n753) );
  XNOR2_X2 U604 ( .A(A[5]), .B(B[4]), .ZN(n755) );
  XNOR2_X2 U606 ( .A(A[5]), .B(B[2]), .ZN(n757) );
  XNOR2_X2 U607 ( .A(A[5]), .B(B[1]), .ZN(n758) );
  XNOR2_X2 U608 ( .A(B[0]), .B(A[5]), .ZN(n759) );
  OR2_X2 U609 ( .A1(B[0]), .A2(n975), .ZN(n760) );
  OAI22_X2 U611 ( .A1(n12), .A2(n974), .B1(n777), .B2(n965), .ZN(n521) );
  OAI22_X2 U614 ( .A1(n12), .A2(n762), .B1(n965), .B2(n761), .ZN(n626) );
  OAI22_X2 U615 ( .A1(n12), .A2(n763), .B1(n965), .B2(n762), .ZN(n627) );
  OAI22_X2 U616 ( .A1(n12), .A2(n764), .B1(n965), .B2(n763), .ZN(n628) );
  OAI22_X2 U617 ( .A1(n12), .A2(n765), .B1(n965), .B2(n764), .ZN(n629) );
  OAI22_X2 U618 ( .A1(n12), .A2(n766), .B1(n965), .B2(n765), .ZN(n630) );
  OAI22_X2 U619 ( .A1(n12), .A2(n767), .B1(n965), .B2(n766), .ZN(n631) );
  OAI22_X2 U620 ( .A1(n12), .A2(n768), .B1(n965), .B2(n767), .ZN(n632) );
  OAI22_X2 U621 ( .A1(n12), .A2(n769), .B1(n965), .B2(n768), .ZN(n633) );
  OAI22_X2 U622 ( .A1(n12), .A2(n770), .B1(n965), .B2(n769), .ZN(n634) );
  OAI22_X2 U623 ( .A1(n12), .A2(n771), .B1(n965), .B2(n770), .ZN(n635) );
  OAI22_X2 U624 ( .A1(n12), .A2(n772), .B1(n965), .B2(n771), .ZN(n636) );
  OAI22_X2 U625 ( .A1(n12), .A2(n773), .B1(n965), .B2(n772), .ZN(n637) );
  OAI22_X2 U626 ( .A1(n12), .A2(n774), .B1(n965), .B2(n773), .ZN(n638) );
  OAI22_X2 U627 ( .A1(n12), .A2(n775), .B1(n965), .B2(n774), .ZN(n639) );
  OAI22_X2 U628 ( .A1(n12), .A2(n776), .B1(n965), .B2(n775), .ZN(n640) );
  AND2_X2 U629 ( .A1(B[0]), .A2(n948), .ZN(n641) );
  XNOR2_X2 U631 ( .A(A[3]), .B(B[15]), .ZN(n761) );
  XNOR2_X2 U632 ( .A(A[3]), .B(B[14]), .ZN(n762) );
  XNOR2_X2 U633 ( .A(A[3]), .B(B[13]), .ZN(n763) );
  XNOR2_X2 U634 ( .A(A[3]), .B(B[12]), .ZN(n764) );
  XNOR2_X2 U635 ( .A(A[3]), .B(B[11]), .ZN(n765) );
  XNOR2_X2 U636 ( .A(A[3]), .B(B[10]), .ZN(n766) );
  XNOR2_X2 U637 ( .A(A[3]), .B(B[9]), .ZN(n767) );
  XNOR2_X2 U638 ( .A(A[3]), .B(B[8]), .ZN(n768) );
  XNOR2_X2 U639 ( .A(A[3]), .B(B[7]), .ZN(n769) );
  XNOR2_X2 U640 ( .A(A[3]), .B(B[6]), .ZN(n770) );
  XNOR2_X2 U641 ( .A(A[3]), .B(B[5]), .ZN(n771) );
  XNOR2_X2 U642 ( .A(A[3]), .B(B[4]), .ZN(n772) );
  XNOR2_X2 U644 ( .A(A[3]), .B(B[2]), .ZN(n774) );
  XNOR2_X2 U645 ( .A(A[3]), .B(B[1]), .ZN(n775) );
  XNOR2_X2 U646 ( .A(B[0]), .B(A[3]), .ZN(n776) );
  OR2_X2 U647 ( .A1(B[0]), .A2(n974), .ZN(n777) );
  OAI22_X2 U649 ( .A1(n6), .A2(n972), .B1(n794), .B2(n834), .ZN(n522) );
  OAI22_X2 U652 ( .A1(n6), .A2(n779), .B1(n778), .B2(n834), .ZN(n643) );
  OAI22_X2 U653 ( .A1(n6), .A2(n780), .B1(n779), .B2(n834), .ZN(n644) );
  OAI22_X2 U654 ( .A1(n6), .A2(n781), .B1(n780), .B2(n834), .ZN(n645) );
  OAI22_X2 U655 ( .A1(n6), .A2(n782), .B1(n781), .B2(n834), .ZN(n646) );
  OAI22_X2 U656 ( .A1(n6), .A2(n783), .B1(n782), .B2(n834), .ZN(n647) );
  OAI22_X2 U657 ( .A1(n6), .A2(n784), .B1(n783), .B2(n834), .ZN(n648) );
  OAI22_X2 U658 ( .A1(n6), .A2(n785), .B1(n784), .B2(n834), .ZN(n649) );
  OAI22_X2 U659 ( .A1(n6), .A2(n786), .B1(n785), .B2(n834), .ZN(n650) );
  OAI22_X2 U660 ( .A1(n6), .A2(n787), .B1(n786), .B2(n834), .ZN(n651) );
  OAI22_X2 U661 ( .A1(n6), .A2(n788), .B1(n787), .B2(n834), .ZN(n652) );
  OAI22_X2 U662 ( .A1(n6), .A2(n789), .B1(n788), .B2(n834), .ZN(n653) );
  OAI22_X2 U663 ( .A1(n6), .A2(n790), .B1(n789), .B2(n834), .ZN(n654) );
  OAI22_X2 U665 ( .A1(n6), .A2(n792), .B1(n791), .B2(n834), .ZN(n656) );
  OAI22_X2 U666 ( .A1(n6), .A2(n793), .B1(n792), .B2(n834), .ZN(n657) );
  AND2_X2 U667 ( .A1(B[0]), .A2(A[0]), .ZN(n658) );
  XNOR2_X2 U669 ( .A(n973), .B(B[15]), .ZN(n778) );
  XNOR2_X2 U670 ( .A(n973), .B(B[14]), .ZN(n779) );
  XNOR2_X2 U671 ( .A(n973), .B(B[13]), .ZN(n780) );
  XNOR2_X2 U672 ( .A(n973), .B(B[12]), .ZN(n781) );
  XNOR2_X2 U673 ( .A(n973), .B(B[11]), .ZN(n782) );
  XNOR2_X2 U674 ( .A(n973), .B(B[10]), .ZN(n783) );
  XNOR2_X2 U675 ( .A(n973), .B(B[9]), .ZN(n784) );
  XNOR2_X2 U676 ( .A(n973), .B(B[8]), .ZN(n785) );
  XNOR2_X2 U677 ( .A(n973), .B(B[7]), .ZN(n786) );
  XNOR2_X2 U678 ( .A(n973), .B(B[6]), .ZN(n787) );
  XNOR2_X2 U679 ( .A(n973), .B(B[5]), .ZN(n788) );
  XNOR2_X2 U680 ( .A(n973), .B(B[4]), .ZN(n789) );
  XNOR2_X2 U682 ( .A(n973), .B(B[2]), .ZN(n791) );
  XNOR2_X2 U683 ( .A(n973), .B(B[1]), .ZN(n792) );
  XNOR2_X2 U684 ( .A(B[0]), .B(n973), .ZN(n793) );
  OR2_X2 U685 ( .A1(B[0]), .A2(n972), .ZN(n794) );
  XOR2_X2 U711 ( .A(A[14]), .B(A[15]), .Z(n811) );
  XOR2_X2 U714 ( .A(A[12]), .B(A[13]), .Z(n812) );
  XOR2_X2 U717 ( .A(A[10]), .B(n979), .Z(n813) );
  XOR2_X2 U720 ( .A(A[8]), .B(A[9]), .Z(n814) );
  XOR2_X2 U723 ( .A(A[6]), .B(A[7]), .Z(n815) );
  XOR2_X2 U726 ( .A(A[4]), .B(A[5]), .Z(n816) );
  XOR2_X2 U729 ( .A(A[2]), .B(A[3]), .Z(n817) );
  XOR2_X2 U732 ( .A(A[0]), .B(n973), .Z(n818) );
  INV_X1 U737 ( .A(A[3]), .ZN(n974) );
  INV_X1 U738 ( .A(A[9]), .ZN(n977) );
  XOR2_X2 U739 ( .A(n238), .B(n243), .Z(n937) );
  XOR2_X2 U740 ( .A(n82), .B(n937), .Z(MAC[26]) );
  NAND2_X2 U741 ( .A1(n238), .A2(n82), .ZN(n938) );
  NAND2_X2 U742 ( .A1(n243), .A2(n82), .ZN(n939) );
  NAND2_X2 U743 ( .A1(n243), .A2(n238), .ZN(n940) );
  NAND3_X2 U744 ( .A1(n940), .A2(n939), .A3(n938), .ZN(n81) );
  XOR2_X2 U745 ( .A(n390), .B(n392), .Z(n941) );
  XOR2_X2 U746 ( .A(n388), .B(n941), .Z(n384) );
  NAND2_X2 U747 ( .A1(n390), .A2(n388), .ZN(n942) );
  NAND2_X2 U748 ( .A1(n392), .A2(n388), .ZN(n943) );
  NAND2_X2 U749 ( .A1(n392), .A2(n390), .ZN(n944) );
  NAND3_X2 U750 ( .A1(n944), .A2(n943), .A3(n942), .ZN(n383) );
  AOI21_X4 U751 ( .B1(n127), .B2(n119), .A(n120), .ZN(n118) );
  XNOR2_X1 U752 ( .A(A[7]), .B(B[8]), .ZN(n734) );
  XNOR2_X1 U753 ( .A(A[7]), .B(B[5]), .ZN(n737) );
  XNOR2_X1 U754 ( .A(A[5]), .B(B[15]), .ZN(n744) );
  XNOR2_X1 U755 ( .A(A[5]), .B(B[5]), .ZN(n754) );
  INV_X1 U756 ( .A(A[5]), .ZN(n975) );
  INV_X1 U757 ( .A(A[13]), .ZN(n980) );
  XOR2_X2 U758 ( .A(A[5]), .B(A[6]), .Z(n945) );
  XOR2_X2 U759 ( .A(A[13]), .B(A[14]), .Z(n946) );
  XOR2_X2 U760 ( .A(n979), .B(A[12]), .Z(n947) );
  XOR2_X2 U761 ( .A(n973), .B(A[2]), .Z(n948) );
  XOR2_X2 U762 ( .A(A[3]), .B(A[4]), .Z(n949) );
  XOR2_X2 U763 ( .A(A[7]), .B(A[8]), .Z(n950) );
  XOR2_X2 U764 ( .A(A[9]), .B(A[10]), .Z(n951) );
  OR2_X4 U765 ( .A1(n658), .A2(C[0]), .ZN(n952) );
  AND2_X4 U766 ( .A1(n952), .A2(n194), .ZN(MAC[0]) );
  XNOR2_X2 U767 ( .A(n51), .B(n77), .ZN(n954) );
  INV_X4 U768 ( .A(n954), .ZN(MAC[31]) );
  XNOR2_X1 U769 ( .A(A[15]), .B(B[3]), .ZN(n671) );
  XNOR2_X1 U770 ( .A(A[5]), .B(B[3]), .ZN(n756) );
  XNOR2_X1 U771 ( .A(n973), .B(B[3]), .ZN(n790) );
  XNOR2_X1 U772 ( .A(A[3]), .B(B[3]), .ZN(n773) );
  XNOR2_X1 U773 ( .A(A[13]), .B(B[3]), .ZN(n688) );
  XNOR2_X1 U774 ( .A(A[7]), .B(B[3]), .ZN(n739) );
  XNOR2_X1 U775 ( .A(n979), .B(B[3]), .ZN(n705) );
  XNOR2_X1 U776 ( .A(A[9]), .B(B[3]), .ZN(n722) );
  AOI21_X2 U777 ( .B1(n115), .B2(n956), .A(n112), .ZN(n110) );
  AOI21_X2 U778 ( .B1(n107), .B2(n957), .A(n104), .ZN(n102) );
  AOI21_X2 U779 ( .B1(n99), .B2(n958), .A(n96), .ZN(n94) );
  AOI21_X2 U780 ( .B1(n91), .B2(n959), .A(n88), .ZN(n86) );
  NAND2_X2 U781 ( .A1(n816), .A2(n966), .ZN(n18) );
  NAND2_X2 U782 ( .A1(n812), .A2(n970), .ZN(n42) );
  INV_X4 U783 ( .A(n945), .ZN(n967) );
  INV_X4 U784 ( .A(n946), .ZN(n971) );
  INV_X4 U785 ( .A(n978), .ZN(n979) );
  INV_X2 U786 ( .A(n145), .ZN(n144) );
  NOR2_X1 U787 ( .A1(n121), .A2(n124), .ZN(n119) );
  INV_X1 U788 ( .A(n148), .ZN(n209) );
  INV_X2 U789 ( .A(n143), .ZN(n141) );
  NOR2_X1 U790 ( .A1(n420), .A2(n431), .ZN(n142) );
  NAND2_X1 U791 ( .A1(n432), .A2(n441), .ZN(n149) );
  OAI22_X1 U792 ( .A1(n778), .A2(n6), .B1(n778), .B2(n834), .ZN(n512) );
  OAI22_X1 U793 ( .A1(n42), .A2(n682), .B1(n970), .B2(n681), .ZN(n546) );
  OAI22_X1 U794 ( .A1(n48), .A2(n665), .B1(n971), .B2(n664), .ZN(n529) );
  OAI21_X1 U795 ( .B1(n126), .B2(n124), .A(n125), .ZN(n123) );
  NAND2_X1 U796 ( .A1(n204), .A2(n122), .ZN(n61) );
  OAI22_X1 U797 ( .A1(n676), .A2(n42), .B1(n676), .B2(n970), .ZN(n494) );
  AOI21_X1 U798 ( .B1(n144), .B2(n135), .A(n136), .ZN(n134) );
  NAND2_X1 U799 ( .A1(n955), .A2(n133), .ZN(n63) );
  NAND2_X1 U800 ( .A1(n208), .A2(n143), .ZN(n65) );
  OAI22_X1 U801 ( .A1(n6), .A2(n791), .B1(n790), .B2(n834), .ZN(n655) );
  OAI21_X2 U802 ( .B1(n121), .B2(n125), .A(n122), .ZN(n120) );
  AOI21_X2 U803 ( .B1(n146), .B2(n154), .A(n147), .ZN(n145) );
  NOR2_X2 U804 ( .A1(n148), .A2(n151), .ZN(n146) );
  OAI21_X2 U805 ( .B1(n148), .B2(n152), .A(n149), .ZN(n147) );
  OAI21_X2 U806 ( .B1(n145), .B2(n128), .A(n129), .ZN(n127) );
  AOI21_X2 U807 ( .B1(n955), .B2(n136), .A(n131), .ZN(n129) );
  OAI21_X2 U808 ( .B1(n118), .B2(n116), .A(n117), .ZN(n115) );
  OAI21_X2 U809 ( .B1(n110), .B2(n108), .A(n109), .ZN(n107) );
  OAI21_X2 U810 ( .B1(n102), .B2(n100), .A(n101), .ZN(n99) );
  OAI21_X2 U811 ( .B1(n94), .B2(n92), .A(n93), .ZN(n91) );
  OAI21_X2 U812 ( .B1(n137), .B2(n143), .A(n138), .ZN(n136) );
  OAI21_X2 U813 ( .B1(n157), .B2(n155), .A(n156), .ZN(n154) );
  NOR2_X2 U814 ( .A1(n137), .A2(n142), .ZN(n135) );
  AOI21_X2 U815 ( .B1(n162), .B2(n963), .A(n159), .ZN(n157) );
  AOI21_X2 U816 ( .B1(n960), .B2(n180), .A(n177), .ZN(n175) );
  OAI21_X2 U817 ( .B1(n163), .B2(n175), .A(n164), .ZN(n162) );
  AOI21_X2 U818 ( .B1(n961), .B2(n171), .A(n166), .ZN(n164) );
  NOR2_X2 U819 ( .A1(n408), .A2(n419), .ZN(n137) );
  NOR2_X2 U820 ( .A1(n364), .A2(n379), .ZN(n121) );
  NOR2_X2 U821 ( .A1(n432), .A2(n441), .ZN(n148) );
  NOR2_X2 U822 ( .A1(n380), .A2(n393), .ZN(n124) );
  NOR2_X2 U823 ( .A1(n442), .A2(n451), .ZN(n151) );
  NOR2_X2 U824 ( .A1(n348), .A2(n363), .ZN(n116) );
  NOR2_X2 U825 ( .A1(n318), .A2(n331), .ZN(n108) );
  NOR2_X2 U826 ( .A1(n452), .A2(n459), .ZN(n155) );
  OR2_X1 U827 ( .A1(n394), .A2(n407), .ZN(n955) );
  OR2_X1 U828 ( .A1(n332), .A2(n347), .ZN(n956) );
  OR2_X1 U829 ( .A1(n304), .A2(n317), .ZN(n957) );
  NOR2_X2 U830 ( .A1(n292), .A2(n303), .ZN(n100) );
  NOR2_X2 U831 ( .A1(n270), .A2(n279), .ZN(n92) );
  OR2_X1 U832 ( .A1(n280), .A2(n291), .ZN(n958) );
  OR2_X1 U833 ( .A1(n260), .A2(n269), .ZN(n959) );
  NOR2_X2 U834 ( .A1(n252), .A2(n259), .ZN(n84) );
  OAI21_X2 U835 ( .B1(n181), .B2(n183), .A(n182), .ZN(n180) );
  OAI21_X2 U836 ( .B1(n86), .B2(n84), .A(n85), .ZN(n83) );
  OR2_X1 U837 ( .A1(n480), .A2(n483), .ZN(n960) );
  OR2_X1 U838 ( .A1(n468), .A2(n473), .ZN(n961) );
  OR2_X1 U839 ( .A1(n474), .A2(n479), .ZN(n962) );
  OR2_X1 U840 ( .A1(n460), .A2(n467), .ZN(n963) );
  AOI21_X2 U841 ( .B1(n964), .B2(n192), .A(n189), .ZN(n187) );
  OAI21_X2 U842 ( .B1(n187), .B2(n185), .A(n186), .ZN(n184) );
  INV_X4 U843 ( .A(n512), .ZN(n642) );
  INV_X4 U844 ( .A(n509), .ZN(n625) );
  NOR2_X2 U845 ( .A1(n484), .A2(n486), .ZN(n181) );
  INV_X4 U846 ( .A(n506), .ZN(n608) );
  NOR2_X2 U847 ( .A1(n488), .A2(n489), .ZN(n185) );
  OR2_X1 U848 ( .A1(n490), .A2(n522), .ZN(n964) );
  INV_X4 U849 ( .A(n503), .ZN(n591) );
  INV_X4 U850 ( .A(n500), .ZN(n574) );
  INV_X4 U851 ( .A(n497), .ZN(n557) );
  INV_X4 U852 ( .A(n494), .ZN(n540) );
  AOI21_X2 U853 ( .B1(n144), .B2(n208), .A(n141), .ZN(n139) );
  AOI21_X2 U854 ( .B1(n174), .B2(n962), .A(n171), .ZN(n169) );
  OAI21_X2 U855 ( .B1(n153), .B2(n151), .A(n152), .ZN(n150) );
  XNOR2_X2 U856 ( .A(C[31]), .B(n221), .ZN(n51) );
  NAND2_X2 U857 ( .A1(n815), .A2(n967), .ZN(n24) );
  NAND2_X2 U858 ( .A1(n814), .A2(n968), .ZN(n30) );
  NAND2_X2 U859 ( .A1(n813), .A2(n969), .ZN(n36) );
  NAND2_X2 U860 ( .A1(n811), .A2(n971), .ZN(n48) );
  NAND2_X2 U861 ( .A1(n817), .A2(n965), .ZN(n12) );
  NAND2_X2 U862 ( .A1(n818), .A2(n834), .ZN(n6) );
  INV_X4 U863 ( .A(A[0]), .ZN(n834) );
  INV_X4 U864 ( .A(A[15]), .ZN(n981) );
  INV_X4 U865 ( .A(A[7]), .ZN(n976) );
  INV_X4 U866 ( .A(n972), .ZN(n973) );
  INV_X4 U867 ( .A(A[1]), .ZN(n972) );
  INV_X4 U868 ( .A(A[11]), .ZN(n978) );
  INV_X4 U869 ( .A(n951), .ZN(n969) );
  INV_X4 U870 ( .A(n948), .ZN(n965) );
  INV_X4 U871 ( .A(n950), .ZN(n968) );
  INV_X4 U872 ( .A(n947), .ZN(n970) );
  INV_X4 U873 ( .A(n949), .ZN(n966) );
  INV_X4 U874 ( .A(n491), .ZN(n523) );
  INV_X4 U875 ( .A(n98), .ZN(n96) );
  INV_X4 U876 ( .A(n90), .ZN(n88) );
  OAI22_X2 U877 ( .A1(n761), .A2(n12), .B1(n761), .B2(n965), .ZN(n509) );
  OAI22_X2 U878 ( .A1(n744), .A2(n18), .B1(n744), .B2(n966), .ZN(n506) );
  OAI22_X2 U879 ( .A1(n727), .A2(n24), .B1(n727), .B2(n967), .ZN(n503) );
  OAI22_X2 U880 ( .A1(n710), .A2(n30), .B1(n710), .B2(n968), .ZN(n500) );
  OAI22_X2 U881 ( .A1(n693), .A2(n36), .B1(n693), .B2(n969), .ZN(n497) );
  OAI22_X2 U882 ( .A1(n659), .A2(n48), .B1(n659), .B2(n971), .ZN(n491) );
  INV_X4 U883 ( .A(C[17]), .ZN(n346) );
  INV_X4 U884 ( .A(C[19]), .ZN(n316) );
  INV_X4 U885 ( .A(C[21]), .ZN(n290) );
  INV_X4 U886 ( .A(C[23]), .ZN(n268) );
  INV_X4 U887 ( .A(C[25]), .ZN(n250) );
  INV_X4 U888 ( .A(C[27]), .ZN(n236) );
  INV_X4 U889 ( .A(C[29]), .ZN(n226) );
  INV_X4 U890 ( .A(n185), .ZN(n217) );
  INV_X4 U891 ( .A(n181), .ZN(n216) );
  INV_X4 U892 ( .A(n155), .ZN(n211) );
  INV_X4 U893 ( .A(n151), .ZN(n210) );
  INV_X4 U894 ( .A(n137), .ZN(n207) );
  INV_X4 U895 ( .A(n124), .ZN(n205) );
  INV_X4 U896 ( .A(n121), .ZN(n204) );
  INV_X4 U897 ( .A(n116), .ZN(n203) );
  INV_X4 U898 ( .A(n108), .ZN(n201) );
  INV_X4 U899 ( .A(n100), .ZN(n199) );
  INV_X4 U900 ( .A(n92), .ZN(n197) );
  INV_X4 U901 ( .A(n84), .ZN(n195) );
  INV_X4 U902 ( .A(n194), .ZN(n192) );
  INV_X4 U903 ( .A(n191), .ZN(n189) );
  INV_X4 U904 ( .A(n184), .ZN(n183) );
  INV_X4 U905 ( .A(n179), .ZN(n177) );
  INV_X4 U906 ( .A(n175), .ZN(n174) );
  INV_X4 U907 ( .A(n173), .ZN(n171) );
  INV_X4 U908 ( .A(n168), .ZN(n166) );
  INV_X4 U909 ( .A(n161), .ZN(n159) );
  INV_X4 U910 ( .A(n154), .ZN(n153) );
  INV_X4 U911 ( .A(n142), .ZN(n208) );
  INV_X4 U912 ( .A(n133), .ZN(n131) );
  INV_X4 U913 ( .A(n127), .ZN(n126) );
  INV_X4 U914 ( .A(n114), .ZN(n112) );
  INV_X4 U915 ( .A(n106), .ZN(n104) );
  XNOR2_X1 U916 ( .A(A[7]), .B(B[7]), .ZN(n735) );
endmodule


module macopertion_3 ( in_a_mac, in_b_mac, bitselect1, clk, min );
  input [15:0] in_a_mac;
  input [15:0] in_b_mac;
  input [3:0] bitselect1;
  output [15:0] min;
  input clk;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18,
         N19, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49,
         N50, N51, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198;
  wire   [31:0] in_c_mac;
  wire   [31:0] out_mac;
  assign min[15] = 1'b0;

  macopertion_3_DW02_mac_1 U1 ( .A({in_a_mac[15:6], n179, in_a_mac[4:0]}), .B(
        {in_b_mac[15:1], n180}), .C(in_c_mac), .TC(1'b1), .MAC(out_mac) );
  DFF_X1 in_c_mac_reg_0_ ( .D(N4), .CK(clk), .Q(in_c_mac[0]) );
  DFF_X1 in_c_mac_reg_1_ ( .D(N5), .CK(clk), .Q(in_c_mac[1]) );
  DFF_X1 in_c_mac_reg_2_ ( .D(N6), .CK(clk), .Q(in_c_mac[2]) );
  DFF_X1 in_c_mac_reg_3_ ( .D(N7), .CK(clk), .Q(in_c_mac[3]) );
  DFF_X1 in_c_mac_reg_4_ ( .D(N8), .CK(clk), .Q(in_c_mac[4]) );
  DFF_X1 in_c_mac_reg_5_ ( .D(N9), .CK(clk), .Q(in_c_mac[5]) );
  DFF_X1 in_c_mac_reg_6_ ( .D(N10), .CK(clk), .Q(in_c_mac[6]) );
  DFF_X1 in_c_mac_reg_7_ ( .D(N11), .CK(clk), .Q(in_c_mac[7]) );
  DFF_X1 in_c_mac_reg_8_ ( .D(N12), .CK(clk), .Q(in_c_mac[8]) );
  DFF_X1 in_c_mac_reg_9_ ( .D(N13), .CK(clk), .Q(in_c_mac[9]) );
  DFF_X1 in_c_mac_reg_10_ ( .D(N14), .CK(clk), .Q(in_c_mac[10]) );
  DFF_X1 in_c_mac_reg_11_ ( .D(N15), .CK(clk), .Q(in_c_mac[11]) );
  DFF_X1 in_c_mac_reg_12_ ( .D(N16), .CK(clk), .Q(in_c_mac[12]) );
  DFF_X1 in_c_mac_reg_13_ ( .D(N17), .CK(clk), .Q(in_c_mac[13]) );
  DFF_X1 in_c_mac_reg_14_ ( .D(N18), .CK(clk), .Q(in_c_mac[14]) );
  DFF_X1 in_c_mac_reg_15_ ( .D(N19), .CK(clk), .Q(in_c_mac[15]) );
  SDFF_X1 in_c_mac_reg_16_ ( .D(out_mac[16]), .SI(1'b0), .SE(n198), .CK(clk), 
        .Q(in_c_mac[16]) );
  SDFF_X1 in_c_mac_reg_17_ ( .D(out_mac[17]), .SI(1'b0), .SE(n198), .CK(clk), 
        .Q(in_c_mac[17]) );
  SDFF_X1 in_c_mac_reg_18_ ( .D(out_mac[18]), .SI(1'b0), .SE(n198), .CK(clk), 
        .Q(in_c_mac[18]) );
  SDFF_X1 in_c_mac_reg_19_ ( .D(out_mac[19]), .SI(1'b0), .SE(n198), .CK(clk), 
        .Q(in_c_mac[19]) );
  SDFF_X1 in_c_mac_reg_20_ ( .D(out_mac[20]), .SI(1'b0), .SE(n198), .CK(clk), 
        .Q(in_c_mac[20]) );
  SDFF_X1 in_c_mac_reg_21_ ( .D(out_mac[21]), .SI(1'b0), .SE(n198), .CK(clk), 
        .Q(in_c_mac[21]) );
  SDFF_X1 in_c_mac_reg_22_ ( .D(out_mac[22]), .SI(1'b0), .SE(n198), .CK(clk), 
        .Q(in_c_mac[22]) );
  SDFF_X1 in_c_mac_reg_23_ ( .D(out_mac[23]), .SI(1'b0), .SE(n198), .CK(clk), 
        .Q(in_c_mac[23]) );
  SDFF_X1 in_c_mac_reg_24_ ( .D(out_mac[24]), .SI(1'b0), .SE(n198), .CK(clk), 
        .Q(in_c_mac[24]) );
  SDFF_X1 in_c_mac_reg_25_ ( .D(out_mac[25]), .SI(1'b0), .SE(n198), .CK(clk), 
        .Q(in_c_mac[25]) );
  SDFF_X1 in_c_mac_reg_26_ ( .D(out_mac[26]), .SI(1'b0), .SE(n198), .CK(clk), 
        .Q(in_c_mac[26]) );
  SDFF_X1 in_c_mac_reg_27_ ( .D(out_mac[27]), .SI(1'b0), .SE(n198), .CK(clk), 
        .Q(in_c_mac[27]) );
  SDFF_X1 in_c_mac_reg_28_ ( .D(out_mac[28]), .SI(1'b0), .SE(n198), .CK(clk), 
        .Q(in_c_mac[28]) );
  SDFF_X1 in_c_mac_reg_29_ ( .D(out_mac[29]), .SI(1'b0), .SE(n198), .CK(clk), 
        .Q(in_c_mac[29]) );
  SDFF_X1 in_c_mac_reg_30_ ( .D(out_mac[30]), .SI(1'b0), .SE(n198), .CK(clk), 
        .Q(in_c_mac[30]) );
  DFF_X1 min_reg_14_ ( .D(N51), .CK(clk), .Q(min[14]) );
  DFF_X1 min_reg_13_ ( .D(N50), .CK(clk), .Q(min[13]) );
  DFF_X1 min_reg_12_ ( .D(N49), .CK(clk), .Q(min[12]) );
  DFF_X1 min_reg_11_ ( .D(N48), .CK(clk), .Q(min[11]) );
  DFF_X1 min_reg_10_ ( .D(N47), .CK(clk), .Q(min[10]) );
  DFF_X1 min_reg_9_ ( .D(N46), .CK(clk), .Q(min[9]) );
  DFF_X1 min_reg_8_ ( .D(N45), .CK(clk), .Q(min[8]) );
  DFF_X1 min_reg_7_ ( .D(N44), .CK(clk), .Q(min[7]) );
  DFF_X1 min_reg_6_ ( .D(N43), .CK(clk), .Q(min[6]) );
  DFF_X1 min_reg_5_ ( .D(N42), .CK(clk), .Q(min[5]) );
  DFF_X1 min_reg_4_ ( .D(N41), .CK(clk), .Q(min[4]) );
  DFF_X1 min_reg_3_ ( .D(N40), .CK(clk), .Q(min[3]) );
  DFF_X1 min_reg_2_ ( .D(N39), .CK(clk), .Q(min[2]) );
  DFF_X1 min_reg_1_ ( .D(N38), .CK(clk), .Q(min[1]) );
  DFF_X1 min_reg_0_ ( .D(N37), .CK(clk), .Q(min[0]) );
  SDFF_X2 in_c_mac_reg_31_ ( .D(out_mac[31]), .SI(1'b0), .SE(n198), .CK(clk), 
        .Q(in_c_mac[31]) );
  BUF_X4 U23 ( .A(in_a_mac[5]), .Z(n179) );
  INV_X4 U24 ( .A(n181), .ZN(n180) );
  INV_X1 U25 ( .A(in_b_mac[0]), .ZN(n181) );
  INV_X4 U26 ( .A(n182), .ZN(n198) );
  OR4_X4 U27 ( .A1(bitselect1[1]), .A2(bitselect1[0]), .A3(bitselect1[3]), 
        .A4(bitselect1[2]), .ZN(n182) );
  AND2_X1 U28 ( .A1(out_mac[15]), .A2(n182), .ZN(N19) );
  AND2_X1 U29 ( .A1(out_mac[14]), .A2(n182), .ZN(N18) );
  AND2_X1 U30 ( .A1(out_mac[13]), .A2(n182), .ZN(N17) );
  AND2_X1 U31 ( .A1(out_mac[12]), .A2(n182), .ZN(N16) );
  AND2_X1 U32 ( .A1(out_mac[11]), .A2(n182), .ZN(N15) );
  AND2_X1 U33 ( .A1(out_mac[10]), .A2(n182), .ZN(N14) );
  AND2_X1 U34 ( .A1(out_mac[9]), .A2(n182), .ZN(N13) );
  AND2_X1 U35 ( .A1(out_mac[8]), .A2(n182), .ZN(N12) );
  AND2_X1 U36 ( .A1(out_mac[7]), .A2(n182), .ZN(N11) );
  AND2_X1 U37 ( .A1(out_mac[6]), .A2(n182), .ZN(N10) );
  AND2_X1 U38 ( .A1(out_mac[5]), .A2(n182), .ZN(N9) );
  AND2_X1 U39 ( .A1(out_mac[4]), .A2(n182), .ZN(N8) );
  AND2_X1 U40 ( .A1(out_mac[3]), .A2(n182), .ZN(N7) );
  AND2_X1 U41 ( .A1(out_mac[2]), .A2(n182), .ZN(N6) );
  AND2_X1 U42 ( .A1(out_mac[1]), .A2(n182), .ZN(N5) );
  AND2_X1 U43 ( .A1(out_mac[0]), .A2(n182), .ZN(N4) );
  INV_X4 U44 ( .A(out_mac[16]), .ZN(n183) );
  NOR2_X2 U45 ( .A1(out_mac[31]), .A2(n183), .ZN(N37) );
  INV_X4 U46 ( .A(out_mac[17]), .ZN(n184) );
  NOR2_X2 U47 ( .A1(out_mac[31]), .A2(n184), .ZN(N38) );
  INV_X4 U48 ( .A(out_mac[18]), .ZN(n185) );
  NOR2_X2 U49 ( .A1(out_mac[31]), .A2(n185), .ZN(N39) );
  INV_X4 U50 ( .A(out_mac[19]), .ZN(n186) );
  NOR2_X2 U51 ( .A1(out_mac[31]), .A2(n186), .ZN(N40) );
  INV_X4 U52 ( .A(out_mac[20]), .ZN(n187) );
  NOR2_X2 U53 ( .A1(out_mac[31]), .A2(n187), .ZN(N41) );
  INV_X4 U54 ( .A(out_mac[21]), .ZN(n188) );
  NOR2_X2 U55 ( .A1(out_mac[31]), .A2(n188), .ZN(N42) );
  INV_X4 U56 ( .A(out_mac[22]), .ZN(n189) );
  NOR2_X2 U57 ( .A1(out_mac[31]), .A2(n189), .ZN(N43) );
  INV_X4 U58 ( .A(out_mac[23]), .ZN(n190) );
  NOR2_X2 U59 ( .A1(out_mac[31]), .A2(n190), .ZN(N44) );
  INV_X4 U60 ( .A(out_mac[24]), .ZN(n191) );
  NOR2_X2 U61 ( .A1(out_mac[31]), .A2(n191), .ZN(N45) );
  INV_X4 U62 ( .A(out_mac[25]), .ZN(n192) );
  NOR2_X2 U63 ( .A1(out_mac[31]), .A2(n192), .ZN(N46) );
  INV_X4 U64 ( .A(out_mac[26]), .ZN(n193) );
  NOR2_X2 U65 ( .A1(out_mac[31]), .A2(n193), .ZN(N47) );
  INV_X4 U66 ( .A(out_mac[27]), .ZN(n194) );
  NOR2_X2 U67 ( .A1(out_mac[31]), .A2(n194), .ZN(N48) );
  INV_X4 U68 ( .A(out_mac[28]), .ZN(n195) );
  NOR2_X2 U69 ( .A1(out_mac[31]), .A2(n195), .ZN(N49) );
  INV_X4 U70 ( .A(out_mac[29]), .ZN(n196) );
  NOR2_X2 U71 ( .A1(out_mac[31]), .A2(n196), .ZN(N50) );
  INV_X4 U72 ( .A(out_mac[30]), .ZN(n197) );
  NOR2_X2 U73 ( .A1(out_mac[31]), .A2(n197), .ZN(N51) );
endmodule


module macopertion_2_DW02_mac_1 ( A, B, C, TC, MAC );
  input [15:0] A;
  input [15:0] B;
  input [31:0] C;
  output [31:0] MAC;
  input TC;
  wire   n6, n12, n18, n24, n28, n30, n36, n42, n48, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n88, n90, n91, n92, n93, n94, n96, n98, n99, n100, n101,
         n102, n104, n106, n107, n108, n109, n110, n112, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n131, n133, n134, n135, n136, n137, n138, n139, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n159, n161, n162, n163, n164, n166,
         n168, n169, n171, n173, n174, n175, n177, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n189, n191, n192, n194, n195, n197,
         n199, n201, n203, n204, n205, n207, n208, n209, n210, n211, n216,
         n217, n221, n222, n223, n224, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n494, n497, n500, n503, n506, n509, n512, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n811, n812, n813, n814, n815, n816, n817, n818, n834,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984;

  FA_X1 U53 ( .A(n223), .B(n222), .CI(n78), .CO(n77), .S(MAC[30]) );
  FA_X1 U54 ( .A(n224), .B(n227), .CI(n79), .CO(n78), .S(MAC[29]) );
  FA_X1 U55 ( .A(n231), .B(n228), .CI(n80), .CO(n79), .S(MAC[28]) );
  FA_X1 U56 ( .A(n237), .B(n232), .CI(n81), .CO(n80), .S(MAC[27]) );
  FA_X1 U57 ( .A(n238), .B(n243), .CI(n82), .CO(n81), .S(MAC[26]) );
  NAND2_X2 U61 ( .A1(n195), .A2(n85), .ZN(n52) );
  NAND2_X2 U64 ( .A1(n252), .A2(n259), .ZN(n85) );
  XNOR2_X2 U65 ( .A(n91), .B(n53), .ZN(MAC[23]) );
  NAND2_X2 U69 ( .A1(n958), .A2(n90), .ZN(n53) );
  NAND2_X2 U72 ( .A1(n260), .A2(n269), .ZN(n90) );
  XOR2_X2 U73 ( .A(n54), .B(n94), .Z(MAC[22]) );
  NAND2_X2 U75 ( .A1(n197), .A2(n93), .ZN(n54) );
  NAND2_X2 U78 ( .A1(n270), .A2(n279), .ZN(n93) );
  XNOR2_X2 U79 ( .A(n99), .B(n55), .ZN(MAC[21]) );
  NAND2_X2 U83 ( .A1(n957), .A2(n98), .ZN(n55) );
  NAND2_X2 U86 ( .A1(n280), .A2(n291), .ZN(n98) );
  XOR2_X2 U87 ( .A(n56), .B(n102), .Z(MAC[20]) );
  NAND2_X2 U89 ( .A1(n199), .A2(n101), .ZN(n56) );
  NAND2_X2 U92 ( .A1(n292), .A2(n303), .ZN(n101) );
  XNOR2_X2 U93 ( .A(n107), .B(n57), .ZN(MAC[19]) );
  NAND2_X2 U97 ( .A1(n956), .A2(n106), .ZN(n57) );
  NAND2_X2 U100 ( .A1(n304), .A2(n317), .ZN(n106) );
  XOR2_X2 U101 ( .A(n58), .B(n110), .Z(MAC[18]) );
  NAND2_X2 U103 ( .A1(n201), .A2(n109), .ZN(n58) );
  NAND2_X2 U106 ( .A1(n318), .A2(n331), .ZN(n109) );
  NAND2_X2 U111 ( .A1(n955), .A2(n114), .ZN(n59) );
  NAND2_X2 U114 ( .A1(n332), .A2(n347), .ZN(n114) );
  NAND2_X2 U117 ( .A1(n203), .A2(n117), .ZN(n60) );
  NAND2_X2 U120 ( .A1(n348), .A2(n363), .ZN(n117) );
  XNOR2_X2 U121 ( .A(n123), .B(n61), .ZN(MAC[15]) );
  NAND2_X2 U128 ( .A1(n364), .A2(n379), .ZN(n122) );
  XOR2_X2 U129 ( .A(n62), .B(n126), .Z(MAC[14]) );
  NAND2_X2 U131 ( .A1(n205), .A2(n125), .ZN(n62) );
  NAND2_X2 U134 ( .A1(n380), .A2(n393), .ZN(n125) );
  XOR2_X2 U135 ( .A(n63), .B(n134), .Z(MAC[13]) );
  NAND2_X2 U138 ( .A1(n954), .A2(n135), .ZN(n128) );
  NAND2_X2 U145 ( .A1(n394), .A2(n407), .ZN(n133) );
  XOR2_X2 U146 ( .A(n64), .B(n139), .Z(MAC[12]) );
  NAND2_X2 U150 ( .A1(n207), .A2(n138), .ZN(n64) );
  NAND2_X2 U153 ( .A1(n408), .A2(n419), .ZN(n138) );
  XNOR2_X2 U154 ( .A(n144), .B(n65), .ZN(MAC[11]) );
  NAND2_X2 U161 ( .A1(n420), .A2(n431), .ZN(n143) );
  XNOR2_X2 U162 ( .A(n150), .B(n66), .ZN(MAC[10]) );
  NAND2_X2 U167 ( .A1(n209), .A2(n149), .ZN(n66) );
  XOR2_X2 U171 ( .A(n67), .B(n153), .Z(MAC[9]) );
  NAND2_X2 U173 ( .A1(n210), .A2(n152), .ZN(n67) );
  NAND2_X2 U176 ( .A1(n442), .A2(n451), .ZN(n152) );
  XOR2_X2 U177 ( .A(n157), .B(n68), .Z(MAC[8]) );
  NAND2_X2 U180 ( .A1(n211), .A2(n156), .ZN(n68) );
  NAND2_X2 U183 ( .A1(n452), .A2(n459), .ZN(n156) );
  XNOR2_X2 U184 ( .A(n69), .B(n162), .ZN(MAC[7]) );
  NAND2_X2 U188 ( .A1(n962), .A2(n161), .ZN(n69) );
  NAND2_X2 U191 ( .A1(n460), .A2(n467), .ZN(n161) );
  XOR2_X2 U192 ( .A(n70), .B(n169), .Z(MAC[6]) );
  NAND2_X2 U194 ( .A1(n960), .A2(n961), .ZN(n163) );
  NAND2_X2 U198 ( .A1(n960), .A2(n168), .ZN(n70) );
  NAND2_X2 U201 ( .A1(n468), .A2(n473), .ZN(n168) );
  XNOR2_X2 U202 ( .A(n174), .B(n71), .ZN(MAC[5]) );
  NAND2_X2 U206 ( .A1(n961), .A2(n173), .ZN(n71) );
  NAND2_X2 U209 ( .A1(n474), .A2(n479), .ZN(n173) );
  XNOR2_X2 U210 ( .A(n72), .B(n180), .ZN(MAC[4]) );
  NAND2_X2 U215 ( .A1(n959), .A2(n179), .ZN(n72) );
  NAND2_X2 U218 ( .A1(n480), .A2(n483), .ZN(n179) );
  XOR2_X2 U219 ( .A(n183), .B(n73), .Z(MAC[3]) );
  NAND2_X2 U221 ( .A1(n216), .A2(n182), .ZN(n73) );
  NAND2_X2 U224 ( .A1(n484), .A2(n486), .ZN(n182) );
  XOR2_X2 U225 ( .A(n187), .B(n74), .Z(MAC[2]) );
  NAND2_X2 U228 ( .A1(n217), .A2(n186), .ZN(n74) );
  NAND2_X2 U231 ( .A1(n488), .A2(n489), .ZN(n186) );
  XNOR2_X2 U232 ( .A(n75), .B(n192), .ZN(MAC[1]) );
  NAND2_X2 U236 ( .A1(n963), .A2(n191), .ZN(n75) );
  NAND2_X2 U239 ( .A1(n490), .A2(n522), .ZN(n191) );
  NAND2_X2 U245 ( .A1(n658), .A2(C[0]), .ZN(n194) );
  FA_X1 U247 ( .A(C[29]), .B(C[30]), .CI(n523), .CO(n221), .S(n222) );
  FA_X1 U248 ( .A(n524), .B(n226), .CI(n229), .CO(n223), .S(n224) );
  FA_X1 U250 ( .A(n233), .B(n540), .CI(n230), .CO(n227), .S(n228) );
  FA_X1 U251 ( .A(C[27]), .B(C[28]), .CI(n525), .CO(n229), .S(n230) );
  FA_X1 U252 ( .A(n234), .B(n241), .CI(n239), .CO(n231), .S(n232) );
  FA_X1 U253 ( .A(n541), .B(n236), .CI(n526), .CO(n233), .S(n234) );
  FA_X1 U255 ( .A(n245), .B(n242), .CI(n240), .CO(n237), .S(n238) );
  FA_X1 U256 ( .A(n557), .B(n527), .CI(n247), .CO(n239), .S(n240) );
  FA_X1 U257 ( .A(C[25]), .B(C[26]), .CI(n542), .CO(n241), .S(n242) );
  FA_X1 U258 ( .A(n246), .B(n248), .CI(n253), .CO(n243), .S(n244) );
  FA_X1 U259 ( .A(n257), .B(n528), .CI(n255), .CO(n245), .S(n246) );
  FA_X1 U260 ( .A(n558), .B(n250), .CI(n543), .CO(n247), .S(n248) );
  FA_X1 U262 ( .A(n254), .B(n263), .CI(n261), .CO(n251), .S(n252) );
  FA_X1 U263 ( .A(n258), .B(n265), .CI(n256), .CO(n253), .S(n254) );
  FA_X1 U264 ( .A(n544), .B(n529), .CI(n574), .CO(n255), .S(n256) );
  FA_X1 U265 ( .A(C[23]), .B(C[24]), .CI(n559), .CO(n257), .S(n258) );
  FA_X1 U266 ( .A(n271), .B(n264), .CI(n262), .CO(n259), .S(n260) );
  FA_X1 U267 ( .A(n266), .B(n275), .CI(n273), .CO(n261), .S(n262) );
  FA_X1 U268 ( .A(n530), .B(n545), .CI(n277), .CO(n263), .S(n264) );
  FA_X1 U269 ( .A(n575), .B(n268), .CI(n560), .CO(n265), .S(n266) );
  FA_X1 U271 ( .A(n281), .B(n274), .CI(n272), .CO(n269), .S(n270) );
  FA_X1 U272 ( .A(n276), .B(n278), .CI(n283), .CO(n271), .S(n272) );
  FA_X1 U273 ( .A(n287), .B(n576), .CI(n285), .CO(n273), .S(n274) );
  FA_X1 U274 ( .A(n531), .B(n546), .CI(n591), .CO(n275), .S(n276) );
  FA_X1 U275 ( .A(C[21]), .B(C[22]), .CI(n561), .CO(n277), .S(n278) );
  FA_X1 U276 ( .A(n293), .B(n284), .CI(n282), .CO(n279), .S(n280) );
  FA_X1 U277 ( .A(n297), .B(n286), .CI(n295), .CO(n281), .S(n282) );
  FA_X1 U278 ( .A(n299), .B(n301), .CI(n288), .CO(n283), .S(n284) );
  FA_X1 U279 ( .A(n547), .B(n532), .CI(n562), .CO(n285), .S(n286) );
  FA_X1 U280 ( .A(n592), .B(n290), .CI(n577), .CO(n287), .S(n288) );
  FA_X1 U282 ( .A(n305), .B(n296), .CI(n294), .CO(n291), .S(n292) );
  FA_X1 U283 ( .A(n298), .B(n309), .CI(n307), .CO(n293), .S(n294) );
  FA_X1 U284 ( .A(n302), .B(n311), .CI(n300), .CO(n295), .S(n296) );
  FA_X1 U285 ( .A(n533), .B(n548), .CI(n313), .CO(n297), .S(n298) );
  FA_X1 U286 ( .A(n593), .B(n563), .CI(n608), .CO(n299), .S(n300) );
  FA_X1 U287 ( .A(C[19]), .B(C[20]), .CI(n578), .CO(n301), .S(n302) );
  FA_X1 U288 ( .A(n319), .B(n308), .CI(n306), .CO(n303), .S(n304) );
  FA_X1 U289 ( .A(n310), .B(n323), .CI(n321), .CO(n305), .S(n306) );
  FA_X1 U290 ( .A(n314), .B(n325), .CI(n312), .CO(n307), .S(n308) );
  FA_X1 U291 ( .A(n329), .B(n549), .CI(n327), .CO(n309), .S(n310) );
  FA_X1 U292 ( .A(n534), .B(n579), .CI(n564), .CO(n311), .S(n312) );
  FA_X1 U293 ( .A(n609), .B(n316), .CI(n594), .CO(n313), .S(n314) );
  FA_X1 U295 ( .A(n333), .B(n322), .CI(n320), .CO(n317), .S(n318) );
  FA_X1 U296 ( .A(n324), .B(n337), .CI(n335), .CO(n319), .S(n320) );
  FA_X1 U297 ( .A(n326), .B(n330), .CI(n328), .CO(n321), .S(n322) );
  FA_X1 U298 ( .A(n341), .B(n343), .CI(n339), .CO(n323), .S(n324) );
  FA_X1 U299 ( .A(n550), .B(n610), .CI(n595), .CO(n325), .S(n326) );
  FA_X1 U300 ( .A(n535), .B(n565), .CI(n625), .CO(n327), .S(n328) );
  FA_X1 U301 ( .A(C[17]), .B(C[18]), .CI(n580), .CO(n329), .S(n330) );
  FA_X1 U302 ( .A(n349), .B(n336), .CI(n334), .CO(n331), .S(n332) );
  FA_X1 U303 ( .A(n338), .B(n353), .CI(n351), .CO(n333), .S(n334) );
  FA_X1 U304 ( .A(n342), .B(n344), .CI(n340), .CO(n335), .S(n336) );
  FA_X1 U305 ( .A(n357), .B(n359), .CI(n355), .CO(n337), .S(n338) );
  FA_X1 U306 ( .A(n566), .B(n581), .CI(n361), .CO(n339), .S(n340) );
  FA_X1 U307 ( .A(n536), .B(n596), .CI(n551), .CO(n341), .S(n342) );
  FA_X1 U308 ( .A(n626), .B(n346), .CI(n611), .CO(n343), .S(n344) );
  FA_X1 U310 ( .A(n365), .B(n352), .CI(n350), .CO(n347), .S(n348) );
  FA_X1 U311 ( .A(n354), .B(n369), .CI(n367), .CO(n349), .S(n350) );
  FA_X1 U312 ( .A(n371), .B(n360), .CI(n356), .CO(n351), .S(n352) );
  FA_X1 U313 ( .A(n373), .B(n375), .CI(n358), .CO(n353), .S(n354) );
  FA_X1 U314 ( .A(n377), .B(n582), .CI(n362), .CO(n355), .S(n356) );
  FA_X1 U315 ( .A(n537), .B(n612), .CI(n552), .CO(n357), .S(n358) );
  FA_X1 U316 ( .A(n627), .B(n567), .CI(n642), .CO(n359), .S(n360) );
  XNOR2_X2 U317 ( .A(n597), .B(C[16]), .ZN(n362) );
  OR2_X2 U318 ( .A1(n597), .A2(C[16]), .ZN(n361) );
  FA_X1 U319 ( .A(n381), .B(n368), .CI(n366), .CO(n363), .S(n364) );
  FA_X1 U320 ( .A(n383), .B(n372), .CI(n370), .CO(n365), .S(n366) );
  FA_X1 U321 ( .A(n376), .B(n374), .CI(n385), .CO(n367), .S(n368) );
  FA_X1 U322 ( .A(n389), .B(n378), .CI(n387), .CO(n369), .S(n370) );
  FA_X1 U323 ( .A(n598), .B(n613), .CI(n391), .CO(n371), .S(n372) );
  FA_X1 U324 ( .A(n553), .B(n568), .CI(n583), .CO(n373), .S(n374) );
  FA_X1 U325 ( .A(n515), .B(n643), .CI(n628), .CO(n375), .S(n376) );
  HA_X1 U326 ( .A(C[15]), .B(n538), .CO(n377), .S(n378) );
  FA_X1 U327 ( .A(n395), .B(n384), .CI(n382), .CO(n379), .S(n380) );
  FA_X1 U328 ( .A(n397), .B(n399), .CI(n386), .CO(n381), .S(n382) );
  FA_X1 U330 ( .A(n403), .B(n405), .CI(n401), .CO(n385), .S(n386) );
  FA_X1 U331 ( .A(n584), .B(n614), .CI(n599), .CO(n387), .S(n388) );
  FA_X1 U332 ( .A(n554), .B(n629), .CI(n569), .CO(n389), .S(n390) );
  FA_X1 U333 ( .A(n539), .B(C[14]), .CI(n644), .CO(n391), .S(n392) );
  FA_X1 U334 ( .A(n398), .B(n409), .CI(n396), .CO(n393), .S(n394) );
  FA_X1 U335 ( .A(n411), .B(n404), .CI(n400), .CO(n395), .S(n396) );
  FA_X1 U336 ( .A(n413), .B(n415), .CI(n402), .CO(n397), .S(n398) );
  FA_X1 U337 ( .A(n417), .B(n615), .CI(n406), .CO(n399), .S(n400) );
  FA_X1 U338 ( .A(n630), .B(n585), .CI(n600), .CO(n401), .S(n402) );
  FA_X1 U339 ( .A(n516), .B(n645), .CI(n570), .CO(n403), .S(n404) );
  HA_X1 U340 ( .A(C[13]), .B(n555), .CO(n405), .S(n406) );
  FA_X1 U341 ( .A(n421), .B(n412), .CI(n410), .CO(n407), .S(n408) );
  FA_X1 U342 ( .A(n414), .B(n416), .CI(n423), .CO(n409), .S(n410) );
  FA_X1 U343 ( .A(n425), .B(n427), .CI(n418), .CO(n411), .S(n412) );
  FA_X1 U344 ( .A(n601), .B(n616), .CI(n429), .CO(n413), .S(n414) );
  FA_X1 U345 ( .A(n571), .B(n631), .CI(n586), .CO(n415), .S(n416) );
  FA_X1 U346 ( .A(n556), .B(C[12]), .CI(n646), .CO(n417), .S(n418) );
  FA_X1 U347 ( .A(n433), .B(n424), .CI(n422), .CO(n419), .S(n420) );
  FA_X1 U348 ( .A(n428), .B(n426), .CI(n435), .CO(n421), .S(n422) );
  FA_X1 U349 ( .A(n430), .B(n439), .CI(n437), .CO(n423), .S(n424) );
  FA_X1 U350 ( .A(n587), .B(n617), .CI(n602), .CO(n425), .S(n426) );
  FA_X1 U351 ( .A(n517), .B(n647), .CI(n632), .CO(n427), .S(n428) );
  HA_X1 U352 ( .A(C[11]), .B(n572), .CO(n429), .S(n430) );
  FA_X1 U353 ( .A(n443), .B(n436), .CI(n434), .CO(n431), .S(n432) );
  FA_X1 U354 ( .A(n438), .B(n440), .CI(n445), .CO(n433), .S(n434) );
  FA_X1 U355 ( .A(n449), .B(n618), .CI(n447), .CO(n435), .S(n436) );
  FA_X1 U356 ( .A(n588), .B(n633), .CI(n603), .CO(n437), .S(n438) );
  FA_X1 U357 ( .A(n573), .B(C[10]), .CI(n648), .CO(n439), .S(n440) );
  FA_X1 U358 ( .A(n453), .B(n446), .CI(n444), .CO(n441), .S(n442) );
  FA_X1 U359 ( .A(n455), .B(n450), .CI(n448), .CO(n443), .S(n444) );
  FA_X1 U360 ( .A(n604), .B(n619), .CI(n457), .CO(n445), .S(n446) );
  FA_X1 U361 ( .A(n518), .B(n649), .CI(n634), .CO(n447), .S(n448) );
  HA_X1 U362 ( .A(C[9]), .B(n589), .CO(n449), .S(n450) );
  FA_X1 U363 ( .A(n461), .B(n456), .CI(n454), .CO(n451), .S(n452) );
  FA_X1 U364 ( .A(n463), .B(n465), .CI(n458), .CO(n453), .S(n454) );
  FA_X1 U365 ( .A(n605), .B(n635), .CI(n620), .CO(n455), .S(n456) );
  FA_X1 U366 ( .A(n590), .B(C[8]), .CI(n650), .CO(n457), .S(n458) );
  FA_X1 U367 ( .A(n464), .B(n469), .CI(n462), .CO(n459), .S(n460) );
  FA_X1 U368 ( .A(n471), .B(n636), .CI(n466), .CO(n461), .S(n462) );
  FA_X1 U369 ( .A(n519), .B(n651), .CI(n621), .CO(n463), .S(n464) );
  HA_X1 U370 ( .A(C[7]), .B(n606), .CO(n465), .S(n466) );
  FA_X1 U371 ( .A(n472), .B(n475), .CI(n470), .CO(n467), .S(n468) );
  FA_X1 U372 ( .A(n622), .B(n637), .CI(n477), .CO(n469), .S(n470) );
  FA_X1 U373 ( .A(n607), .B(C[6]), .CI(n652), .CO(n471), .S(n472) );
  FA_X1 U374 ( .A(n478), .B(n481), .CI(n476), .CO(n473), .S(n474) );
  FA_X1 U375 ( .A(n520), .B(n653), .CI(n638), .CO(n475), .S(n476) );
  HA_X1 U376 ( .A(C[5]), .B(n623), .CO(n477), .S(n478) );
  FA_X1 U377 ( .A(n485), .B(n639), .CI(n482), .CO(n479), .S(n480) );
  FA_X1 U378 ( .A(n624), .B(C[4]), .CI(n654), .CO(n481), .S(n482) );
  FA_X1 U379 ( .A(n521), .B(n640), .CI(n487), .CO(n483), .S(n484) );
  HA_X1 U380 ( .A(C[3]), .B(n655), .CO(n485), .S(n486) );
  FA_X1 U381 ( .A(n641), .B(C[2]), .CI(n656), .CO(n487), .S(n488) );
  HA_X1 U382 ( .A(C[1]), .B(n657), .CO(n489), .S(n490) );
  OAI22_X2 U383 ( .A1(n48), .A2(n984), .B1(n675), .B2(n970), .ZN(n515) );
  OAI22_X2 U386 ( .A1(n48), .A2(n660), .B1(n970), .B2(n659), .ZN(n524) );
  OAI22_X2 U387 ( .A1(n48), .A2(n661), .B1(n970), .B2(n660), .ZN(n525) );
  OAI22_X2 U388 ( .A1(n48), .A2(n662), .B1(n970), .B2(n661), .ZN(n526) );
  OAI22_X2 U389 ( .A1(n48), .A2(n663), .B1(n970), .B2(n662), .ZN(n527) );
  OAI22_X2 U390 ( .A1(n48), .A2(n664), .B1(n970), .B2(n663), .ZN(n528) );
  OAI22_X2 U392 ( .A1(n48), .A2(n666), .B1(n970), .B2(n665), .ZN(n530) );
  OAI22_X2 U393 ( .A1(n48), .A2(n667), .B1(n970), .B2(n666), .ZN(n531) );
  OAI22_X2 U394 ( .A1(n48), .A2(n668), .B1(n970), .B2(n667), .ZN(n532) );
  OAI22_X2 U395 ( .A1(n48), .A2(n669), .B1(n970), .B2(n668), .ZN(n533) );
  OAI22_X2 U396 ( .A1(n48), .A2(n670), .B1(n970), .B2(n669), .ZN(n534) );
  OAI22_X2 U397 ( .A1(n48), .A2(n671), .B1(n970), .B2(n670), .ZN(n535) );
  OAI22_X2 U398 ( .A1(n48), .A2(n672), .B1(n970), .B2(n671), .ZN(n536) );
  OAI22_X2 U399 ( .A1(n48), .A2(n673), .B1(n970), .B2(n672), .ZN(n537) );
  OAI22_X2 U400 ( .A1(n48), .A2(n674), .B1(n970), .B2(n673), .ZN(n538) );
  AND2_X2 U401 ( .A1(B[0]), .A2(n949), .ZN(n539) );
  XNOR2_X2 U403 ( .A(A[15]), .B(B[15]), .ZN(n659) );
  XNOR2_X2 U404 ( .A(A[15]), .B(B[14]), .ZN(n660) );
  XNOR2_X2 U405 ( .A(A[15]), .B(B[13]), .ZN(n661) );
  XNOR2_X2 U406 ( .A(A[15]), .B(B[12]), .ZN(n662) );
  XNOR2_X2 U407 ( .A(A[15]), .B(B[11]), .ZN(n663) );
  XNOR2_X2 U408 ( .A(A[15]), .B(B[10]), .ZN(n664) );
  XNOR2_X2 U409 ( .A(A[15]), .B(B[9]), .ZN(n665) );
  XNOR2_X2 U410 ( .A(A[15]), .B(B[8]), .ZN(n666) );
  XNOR2_X2 U411 ( .A(A[15]), .B(B[7]), .ZN(n667) );
  XNOR2_X2 U412 ( .A(A[15]), .B(B[6]), .ZN(n668) );
  XNOR2_X2 U413 ( .A(A[15]), .B(B[5]), .ZN(n669) );
  XNOR2_X2 U414 ( .A(A[15]), .B(B[4]), .ZN(n670) );
  XNOR2_X2 U416 ( .A(A[15]), .B(B[2]), .ZN(n672) );
  XNOR2_X2 U417 ( .A(A[15]), .B(B[1]), .ZN(n673) );
  XNOR2_X2 U418 ( .A(B[0]), .B(A[15]), .ZN(n674) );
  OR2_X2 U419 ( .A1(B[0]), .A2(n984), .ZN(n675) );
  OAI22_X2 U421 ( .A1(n42), .A2(n983), .B1(n692), .B2(n969), .ZN(n516) );
  OAI22_X2 U424 ( .A1(n42), .A2(n677), .B1(n969), .B2(n676), .ZN(n541) );
  OAI22_X2 U425 ( .A1(n42), .A2(n678), .B1(n969), .B2(n677), .ZN(n542) );
  OAI22_X2 U426 ( .A1(n42), .A2(n679), .B1(n969), .B2(n678), .ZN(n543) );
  OAI22_X2 U427 ( .A1(n42), .A2(n680), .B1(n969), .B2(n679), .ZN(n544) );
  OAI22_X2 U428 ( .A1(n42), .A2(n681), .B1(n969), .B2(n680), .ZN(n545) );
  OAI22_X2 U430 ( .A1(n42), .A2(n683), .B1(n969), .B2(n682), .ZN(n547) );
  OAI22_X2 U431 ( .A1(n42), .A2(n684), .B1(n969), .B2(n683), .ZN(n548) );
  OAI22_X2 U432 ( .A1(n42), .A2(n685), .B1(n969), .B2(n684), .ZN(n549) );
  OAI22_X2 U433 ( .A1(n42), .A2(n686), .B1(n969), .B2(n685), .ZN(n550) );
  OAI22_X2 U434 ( .A1(n42), .A2(n687), .B1(n969), .B2(n686), .ZN(n551) );
  OAI22_X2 U435 ( .A1(n42), .A2(n688), .B1(n969), .B2(n687), .ZN(n552) );
  OAI22_X2 U436 ( .A1(n42), .A2(n689), .B1(n969), .B2(n688), .ZN(n553) );
  OAI22_X2 U437 ( .A1(n42), .A2(n690), .B1(n969), .B2(n689), .ZN(n554) );
  OAI22_X2 U438 ( .A1(n42), .A2(n691), .B1(n969), .B2(n690), .ZN(n555) );
  AND2_X2 U439 ( .A1(B[0]), .A2(n950), .ZN(n556) );
  XNOR2_X2 U441 ( .A(A[13]), .B(B[15]), .ZN(n676) );
  XNOR2_X2 U442 ( .A(A[13]), .B(B[14]), .ZN(n677) );
  XNOR2_X2 U443 ( .A(A[13]), .B(B[13]), .ZN(n678) );
  XNOR2_X2 U444 ( .A(A[13]), .B(B[12]), .ZN(n679) );
  XNOR2_X2 U445 ( .A(A[13]), .B(B[11]), .ZN(n680) );
  XNOR2_X2 U446 ( .A(A[13]), .B(B[10]), .ZN(n681) );
  XNOR2_X2 U447 ( .A(A[13]), .B(B[9]), .ZN(n682) );
  XNOR2_X2 U448 ( .A(A[13]), .B(B[8]), .ZN(n683) );
  XNOR2_X2 U449 ( .A(A[13]), .B(B[7]), .ZN(n684) );
  XNOR2_X2 U450 ( .A(A[13]), .B(B[6]), .ZN(n685) );
  XNOR2_X2 U451 ( .A(A[13]), .B(B[5]), .ZN(n686) );
  XNOR2_X2 U452 ( .A(A[13]), .B(B[4]), .ZN(n687) );
  XNOR2_X2 U454 ( .A(A[13]), .B(B[2]), .ZN(n689) );
  XNOR2_X2 U455 ( .A(A[13]), .B(B[1]), .ZN(n690) );
  XNOR2_X2 U456 ( .A(B[0]), .B(A[13]), .ZN(n691) );
  OR2_X2 U457 ( .A1(B[0]), .A2(n983), .ZN(n692) );
  OAI22_X2 U459 ( .A1(n36), .A2(n981), .B1(n709), .B2(n968), .ZN(n517) );
  OAI22_X2 U462 ( .A1(n36), .A2(n694), .B1(n968), .B2(n693), .ZN(n558) );
  OAI22_X2 U463 ( .A1(n36), .A2(n695), .B1(n968), .B2(n694), .ZN(n559) );
  OAI22_X2 U464 ( .A1(n36), .A2(n696), .B1(n968), .B2(n695), .ZN(n560) );
  OAI22_X2 U465 ( .A1(n36), .A2(n697), .B1(n968), .B2(n696), .ZN(n561) );
  OAI22_X2 U466 ( .A1(n36), .A2(n698), .B1(n968), .B2(n697), .ZN(n562) );
  OAI22_X2 U467 ( .A1(n36), .A2(n699), .B1(n968), .B2(n698), .ZN(n563) );
  OAI22_X2 U468 ( .A1(n36), .A2(n700), .B1(n968), .B2(n699), .ZN(n564) );
  OAI22_X2 U469 ( .A1(n36), .A2(n701), .B1(n968), .B2(n700), .ZN(n565) );
  OAI22_X2 U470 ( .A1(n36), .A2(n702), .B1(n968), .B2(n701), .ZN(n566) );
  OAI22_X2 U471 ( .A1(n36), .A2(n703), .B1(n968), .B2(n702), .ZN(n567) );
  OAI22_X2 U472 ( .A1(n36), .A2(n704), .B1(n968), .B2(n703), .ZN(n568) );
  OAI22_X2 U473 ( .A1(n36), .A2(n705), .B1(n968), .B2(n704), .ZN(n569) );
  OAI22_X2 U474 ( .A1(n36), .A2(n706), .B1(n968), .B2(n705), .ZN(n570) );
  OAI22_X2 U475 ( .A1(n36), .A2(n707), .B1(n968), .B2(n706), .ZN(n571) );
  OAI22_X2 U476 ( .A1(n36), .A2(n708), .B1(n968), .B2(n707), .ZN(n572) );
  AND2_X2 U477 ( .A1(B[0]), .A2(n948), .ZN(n573) );
  XNOR2_X2 U479 ( .A(n982), .B(B[15]), .ZN(n693) );
  XNOR2_X2 U480 ( .A(n982), .B(B[14]), .ZN(n694) );
  XNOR2_X2 U481 ( .A(n982), .B(B[13]), .ZN(n695) );
  XNOR2_X2 U482 ( .A(n982), .B(B[12]), .ZN(n696) );
  XNOR2_X2 U483 ( .A(n982), .B(B[11]), .ZN(n697) );
  XNOR2_X2 U484 ( .A(n982), .B(B[10]), .ZN(n698) );
  XNOR2_X2 U485 ( .A(n982), .B(B[9]), .ZN(n699) );
  XNOR2_X2 U486 ( .A(n982), .B(B[8]), .ZN(n700) );
  XNOR2_X2 U487 ( .A(n982), .B(B[7]), .ZN(n701) );
  XNOR2_X2 U488 ( .A(n982), .B(B[6]), .ZN(n702) );
  XNOR2_X2 U489 ( .A(n982), .B(B[5]), .ZN(n703) );
  XNOR2_X2 U490 ( .A(n982), .B(B[4]), .ZN(n704) );
  XNOR2_X2 U492 ( .A(n982), .B(B[2]), .ZN(n706) );
  XNOR2_X2 U493 ( .A(n982), .B(B[1]), .ZN(n707) );
  XNOR2_X2 U494 ( .A(B[0]), .B(n982), .ZN(n708) );
  OR2_X2 U495 ( .A1(B[0]), .A2(n981), .ZN(n709) );
  OAI22_X2 U497 ( .A1(n30), .A2(n979), .B1(n726), .B2(n28), .ZN(n518) );
  OAI22_X2 U500 ( .A1(n30), .A2(n711), .B1(n28), .B2(n710), .ZN(n575) );
  OAI22_X2 U501 ( .A1(n30), .A2(n712), .B1(n28), .B2(n711), .ZN(n576) );
  OAI22_X2 U502 ( .A1(n30), .A2(n713), .B1(n28), .B2(n712), .ZN(n577) );
  OAI22_X2 U503 ( .A1(n30), .A2(n714), .B1(n28), .B2(n713), .ZN(n578) );
  OAI22_X2 U504 ( .A1(n30), .A2(n715), .B1(n28), .B2(n714), .ZN(n579) );
  OAI22_X2 U505 ( .A1(n30), .A2(n716), .B1(n28), .B2(n715), .ZN(n580) );
  OAI22_X2 U506 ( .A1(n30), .A2(n717), .B1(n28), .B2(n716), .ZN(n581) );
  OAI22_X2 U507 ( .A1(n30), .A2(n718), .B1(n28), .B2(n717), .ZN(n582) );
  OAI22_X2 U508 ( .A1(n30), .A2(n719), .B1(n28), .B2(n718), .ZN(n583) );
  OAI22_X2 U509 ( .A1(n30), .A2(n720), .B1(n28), .B2(n719), .ZN(n584) );
  OAI22_X2 U510 ( .A1(n30), .A2(n721), .B1(n28), .B2(n720), .ZN(n585) );
  OAI22_X2 U511 ( .A1(n30), .A2(n722), .B1(n28), .B2(n721), .ZN(n586) );
  OAI22_X2 U512 ( .A1(n30), .A2(n723), .B1(n28), .B2(n722), .ZN(n587) );
  OAI22_X2 U513 ( .A1(n30), .A2(n724), .B1(n28), .B2(n723), .ZN(n588) );
  OAI22_X2 U514 ( .A1(n30), .A2(n725), .B1(n28), .B2(n724), .ZN(n589) );
  AND2_X2 U515 ( .A1(B[0]), .A2(n967), .ZN(n590) );
  XNOR2_X2 U517 ( .A(n980), .B(B[15]), .ZN(n710) );
  XNOR2_X2 U518 ( .A(n980), .B(B[14]), .ZN(n711) );
  XNOR2_X2 U519 ( .A(n980), .B(B[13]), .ZN(n712) );
  XNOR2_X2 U520 ( .A(n980), .B(B[12]), .ZN(n713) );
  XNOR2_X2 U521 ( .A(n980), .B(B[11]), .ZN(n714) );
  XNOR2_X2 U522 ( .A(n980), .B(B[10]), .ZN(n715) );
  XNOR2_X2 U523 ( .A(n980), .B(B[9]), .ZN(n716) );
  XNOR2_X2 U524 ( .A(n980), .B(B[8]), .ZN(n717) );
  XNOR2_X2 U525 ( .A(n980), .B(B[7]), .ZN(n718) );
  XNOR2_X2 U526 ( .A(n980), .B(B[6]), .ZN(n719) );
  XNOR2_X2 U527 ( .A(n980), .B(B[5]), .ZN(n720) );
  XNOR2_X2 U528 ( .A(n980), .B(B[4]), .ZN(n721) );
  XNOR2_X2 U530 ( .A(n980), .B(B[2]), .ZN(n723) );
  XNOR2_X2 U531 ( .A(n980), .B(B[1]), .ZN(n724) );
  XNOR2_X2 U532 ( .A(B[0]), .B(n980), .ZN(n725) );
  OR2_X2 U533 ( .A1(B[0]), .A2(n979), .ZN(n726) );
  OAI22_X2 U535 ( .A1(n24), .A2(n977), .B1(n743), .B2(n966), .ZN(n519) );
  OAI22_X2 U538 ( .A1(n24), .A2(n728), .B1(n966), .B2(n727), .ZN(n592) );
  OAI22_X2 U539 ( .A1(n24), .A2(n729), .B1(n966), .B2(n728), .ZN(n593) );
  OAI22_X2 U540 ( .A1(n24), .A2(n730), .B1(n966), .B2(n729), .ZN(n594) );
  OAI22_X2 U541 ( .A1(n24), .A2(n731), .B1(n966), .B2(n730), .ZN(n595) );
  OAI22_X2 U542 ( .A1(n24), .A2(n732), .B1(n966), .B2(n731), .ZN(n596) );
  OAI22_X2 U543 ( .A1(n24), .A2(n733), .B1(n966), .B2(n732), .ZN(n597) );
  OAI22_X2 U544 ( .A1(n24), .A2(n734), .B1(n966), .B2(n733), .ZN(n598) );
  OAI22_X2 U545 ( .A1(n24), .A2(n735), .B1(n966), .B2(n734), .ZN(n599) );
  OAI22_X2 U546 ( .A1(n24), .A2(n736), .B1(n966), .B2(n735), .ZN(n600) );
  OAI22_X2 U547 ( .A1(n24), .A2(n737), .B1(n966), .B2(n736), .ZN(n601) );
  OAI22_X2 U548 ( .A1(n24), .A2(n738), .B1(n966), .B2(n737), .ZN(n602) );
  OAI22_X2 U549 ( .A1(n24), .A2(n739), .B1(n966), .B2(n738), .ZN(n603) );
  OAI22_X2 U550 ( .A1(n24), .A2(n740), .B1(n966), .B2(n739), .ZN(n604) );
  OAI22_X2 U551 ( .A1(n24), .A2(n741), .B1(n966), .B2(n740), .ZN(n605) );
  OAI22_X2 U552 ( .A1(n24), .A2(n742), .B1(n966), .B2(n741), .ZN(n606) );
  AND2_X2 U553 ( .A1(B[0]), .A2(n947), .ZN(n607) );
  XNOR2_X2 U555 ( .A(n978), .B(B[15]), .ZN(n727) );
  XNOR2_X2 U556 ( .A(n978), .B(B[14]), .ZN(n728) );
  XNOR2_X2 U557 ( .A(n978), .B(B[13]), .ZN(n729) );
  XNOR2_X2 U558 ( .A(n978), .B(B[12]), .ZN(n730) );
  XNOR2_X2 U559 ( .A(n978), .B(B[11]), .ZN(n731) );
  XNOR2_X2 U560 ( .A(n978), .B(B[10]), .ZN(n732) );
  XNOR2_X2 U561 ( .A(n978), .B(B[9]), .ZN(n733) );
  XNOR2_X2 U563 ( .A(n978), .B(B[7]), .ZN(n735) );
  XNOR2_X2 U564 ( .A(n978), .B(B[6]), .ZN(n736) );
  XNOR2_X2 U566 ( .A(n978), .B(B[4]), .ZN(n738) );
  XNOR2_X2 U568 ( .A(n978), .B(B[2]), .ZN(n740) );
  XNOR2_X2 U569 ( .A(n978), .B(B[1]), .ZN(n741) );
  XNOR2_X2 U570 ( .A(B[0]), .B(n978), .ZN(n742) );
  OR2_X2 U571 ( .A1(B[0]), .A2(n977), .ZN(n743) );
  OAI22_X2 U573 ( .A1(n18), .A2(n975), .B1(n760), .B2(n965), .ZN(n520) );
  OAI22_X2 U576 ( .A1(n18), .A2(n745), .B1(n965), .B2(n744), .ZN(n609) );
  OAI22_X2 U577 ( .A1(n18), .A2(n746), .B1(n965), .B2(n745), .ZN(n610) );
  OAI22_X2 U578 ( .A1(n18), .A2(n747), .B1(n965), .B2(n746), .ZN(n611) );
  OAI22_X2 U579 ( .A1(n18), .A2(n748), .B1(n965), .B2(n747), .ZN(n612) );
  OAI22_X2 U580 ( .A1(n18), .A2(n749), .B1(n965), .B2(n748), .ZN(n613) );
  OAI22_X2 U581 ( .A1(n18), .A2(n750), .B1(n965), .B2(n749), .ZN(n614) );
  OAI22_X2 U582 ( .A1(n18), .A2(n751), .B1(n965), .B2(n750), .ZN(n615) );
  OAI22_X2 U583 ( .A1(n18), .A2(n752), .B1(n965), .B2(n751), .ZN(n616) );
  OAI22_X2 U584 ( .A1(n18), .A2(n753), .B1(n965), .B2(n752), .ZN(n617) );
  OAI22_X2 U585 ( .A1(n18), .A2(n754), .B1(n965), .B2(n753), .ZN(n618) );
  OAI22_X2 U586 ( .A1(n18), .A2(n755), .B1(n965), .B2(n754), .ZN(n619) );
  OAI22_X2 U587 ( .A1(n18), .A2(n756), .B1(n965), .B2(n755), .ZN(n620) );
  OAI22_X2 U588 ( .A1(n18), .A2(n757), .B1(n965), .B2(n756), .ZN(n621) );
  OAI22_X2 U589 ( .A1(n18), .A2(n758), .B1(n965), .B2(n757), .ZN(n622) );
  OAI22_X2 U590 ( .A1(n18), .A2(n759), .B1(n965), .B2(n758), .ZN(n623) );
  AND2_X2 U591 ( .A1(B[0]), .A2(n946), .ZN(n624) );
  XNOR2_X2 U593 ( .A(n976), .B(B[15]), .ZN(n744) );
  XNOR2_X2 U594 ( .A(n976), .B(B[14]), .ZN(n745) );
  XNOR2_X2 U595 ( .A(n976), .B(B[13]), .ZN(n746) );
  XNOR2_X2 U596 ( .A(n976), .B(B[12]), .ZN(n747) );
  XNOR2_X2 U597 ( .A(n976), .B(B[11]), .ZN(n748) );
  XNOR2_X2 U598 ( .A(n976), .B(B[10]), .ZN(n749) );
  XNOR2_X2 U599 ( .A(n976), .B(B[9]), .ZN(n750) );
  XNOR2_X2 U600 ( .A(n976), .B(B[8]), .ZN(n751) );
  XNOR2_X2 U601 ( .A(n976), .B(B[7]), .ZN(n752) );
  XNOR2_X2 U602 ( .A(n976), .B(B[6]), .ZN(n753) );
  XNOR2_X2 U603 ( .A(n976), .B(B[5]), .ZN(n754) );
  XNOR2_X2 U604 ( .A(n976), .B(B[4]), .ZN(n755) );
  XNOR2_X2 U606 ( .A(n976), .B(B[2]), .ZN(n757) );
  XNOR2_X2 U607 ( .A(n976), .B(B[1]), .ZN(n758) );
  XNOR2_X2 U608 ( .A(B[0]), .B(n976), .ZN(n759) );
  OR2_X2 U609 ( .A1(B[0]), .A2(n975), .ZN(n760) );
  OAI22_X2 U611 ( .A1(n12), .A2(n973), .B1(n777), .B2(n964), .ZN(n521) );
  OAI22_X2 U614 ( .A1(n12), .A2(n762), .B1(n964), .B2(n761), .ZN(n626) );
  OAI22_X2 U615 ( .A1(n12), .A2(n763), .B1(n964), .B2(n762), .ZN(n627) );
  OAI22_X2 U616 ( .A1(n12), .A2(n764), .B1(n964), .B2(n763), .ZN(n628) );
  OAI22_X2 U617 ( .A1(n12), .A2(n765), .B1(n964), .B2(n764), .ZN(n629) );
  OAI22_X2 U618 ( .A1(n12), .A2(n766), .B1(n964), .B2(n765), .ZN(n630) );
  OAI22_X2 U619 ( .A1(n12), .A2(n767), .B1(n964), .B2(n766), .ZN(n631) );
  OAI22_X2 U620 ( .A1(n12), .A2(n768), .B1(n964), .B2(n767), .ZN(n632) );
  OAI22_X2 U621 ( .A1(n12), .A2(n769), .B1(n964), .B2(n768), .ZN(n633) );
  OAI22_X2 U622 ( .A1(n12), .A2(n770), .B1(n964), .B2(n769), .ZN(n634) );
  OAI22_X2 U623 ( .A1(n12), .A2(n771), .B1(n964), .B2(n770), .ZN(n635) );
  OAI22_X2 U624 ( .A1(n12), .A2(n772), .B1(n964), .B2(n771), .ZN(n636) );
  OAI22_X2 U625 ( .A1(n12), .A2(n773), .B1(n964), .B2(n772), .ZN(n637) );
  OAI22_X2 U626 ( .A1(n12), .A2(n774), .B1(n964), .B2(n773), .ZN(n638) );
  OAI22_X2 U627 ( .A1(n12), .A2(n775), .B1(n964), .B2(n774), .ZN(n639) );
  OAI22_X2 U628 ( .A1(n12), .A2(n776), .B1(n964), .B2(n775), .ZN(n640) );
  AND2_X2 U629 ( .A1(B[0]), .A2(n945), .ZN(n641) );
  XNOR2_X2 U631 ( .A(n974), .B(B[15]), .ZN(n761) );
  XNOR2_X2 U632 ( .A(n974), .B(B[14]), .ZN(n762) );
  XNOR2_X2 U633 ( .A(n974), .B(B[13]), .ZN(n763) );
  XNOR2_X2 U634 ( .A(n974), .B(B[12]), .ZN(n764) );
  XNOR2_X2 U635 ( .A(n974), .B(B[11]), .ZN(n765) );
  XNOR2_X2 U636 ( .A(n974), .B(B[10]), .ZN(n766) );
  XNOR2_X2 U637 ( .A(n974), .B(B[9]), .ZN(n767) );
  XNOR2_X2 U638 ( .A(n974), .B(B[8]), .ZN(n768) );
  XNOR2_X2 U639 ( .A(n974), .B(B[7]), .ZN(n769) );
  XNOR2_X2 U640 ( .A(n974), .B(B[6]), .ZN(n770) );
  XNOR2_X2 U641 ( .A(n974), .B(B[5]), .ZN(n771) );
  XNOR2_X2 U642 ( .A(n974), .B(B[4]), .ZN(n772) );
  XNOR2_X2 U644 ( .A(n974), .B(B[2]), .ZN(n774) );
  XNOR2_X2 U645 ( .A(n974), .B(B[1]), .ZN(n775) );
  XNOR2_X2 U646 ( .A(B[0]), .B(n974), .ZN(n776) );
  OR2_X2 U647 ( .A1(B[0]), .A2(n973), .ZN(n777) );
  OAI22_X2 U649 ( .A1(n6), .A2(n971), .B1(n794), .B2(n834), .ZN(n522) );
  OAI22_X2 U652 ( .A1(n6), .A2(n779), .B1(n778), .B2(n834), .ZN(n643) );
  OAI22_X2 U653 ( .A1(n6), .A2(n780), .B1(n779), .B2(n834), .ZN(n644) );
  OAI22_X2 U654 ( .A1(n6), .A2(n781), .B1(n780), .B2(n834), .ZN(n645) );
  OAI22_X2 U655 ( .A1(n6), .A2(n782), .B1(n781), .B2(n834), .ZN(n646) );
  OAI22_X2 U656 ( .A1(n6), .A2(n783), .B1(n782), .B2(n834), .ZN(n647) );
  OAI22_X2 U657 ( .A1(n6), .A2(n784), .B1(n783), .B2(n834), .ZN(n648) );
  OAI22_X2 U658 ( .A1(n6), .A2(n785), .B1(n784), .B2(n834), .ZN(n649) );
  OAI22_X2 U659 ( .A1(n6), .A2(n786), .B1(n785), .B2(n834), .ZN(n650) );
  OAI22_X2 U660 ( .A1(n6), .A2(n787), .B1(n786), .B2(n834), .ZN(n651) );
  OAI22_X2 U661 ( .A1(n6), .A2(n788), .B1(n787), .B2(n834), .ZN(n652) );
  OAI22_X2 U662 ( .A1(n6), .A2(n789), .B1(n788), .B2(n834), .ZN(n653) );
  OAI22_X2 U663 ( .A1(n6), .A2(n790), .B1(n789), .B2(n834), .ZN(n654) );
  OAI22_X2 U665 ( .A1(n6), .A2(n792), .B1(n791), .B2(n834), .ZN(n656) );
  OAI22_X2 U666 ( .A1(n6), .A2(n793), .B1(n792), .B2(n834), .ZN(n657) );
  AND2_X2 U667 ( .A1(B[0]), .A2(A[0]), .ZN(n658) );
  XNOR2_X2 U669 ( .A(n972), .B(B[15]), .ZN(n778) );
  XNOR2_X2 U670 ( .A(n972), .B(B[14]), .ZN(n779) );
  XNOR2_X2 U671 ( .A(n972), .B(B[13]), .ZN(n780) );
  XNOR2_X2 U672 ( .A(n972), .B(B[12]), .ZN(n781) );
  XNOR2_X2 U673 ( .A(n972), .B(B[11]), .ZN(n782) );
  XNOR2_X2 U674 ( .A(n972), .B(B[10]), .ZN(n783) );
  XNOR2_X2 U675 ( .A(n972), .B(B[9]), .ZN(n784) );
  XNOR2_X2 U676 ( .A(n972), .B(B[8]), .ZN(n785) );
  XNOR2_X2 U677 ( .A(n972), .B(B[7]), .ZN(n786) );
  XNOR2_X2 U678 ( .A(n972), .B(B[6]), .ZN(n787) );
  XNOR2_X2 U679 ( .A(n972), .B(B[5]), .ZN(n788) );
  XNOR2_X2 U680 ( .A(n972), .B(B[4]), .ZN(n789) );
  XNOR2_X2 U682 ( .A(n972), .B(B[2]), .ZN(n791) );
  XNOR2_X2 U683 ( .A(n972), .B(B[1]), .ZN(n792) );
  XNOR2_X2 U684 ( .A(B[0]), .B(n972), .ZN(n793) );
  OR2_X2 U685 ( .A1(B[0]), .A2(n971), .ZN(n794) );
  XOR2_X2 U711 ( .A(A[14]), .B(A[15]), .Z(n811) );
  XOR2_X2 U714 ( .A(A[12]), .B(A[13]), .Z(n812) );
  XOR2_X2 U717 ( .A(A[10]), .B(n982), .Z(n813) );
  XOR2_X2 U720 ( .A(A[8]), .B(n980), .Z(n814) );
  XNOR2_X2 U721 ( .A(n978), .B(A[8]), .ZN(n28) );
  XOR2_X2 U723 ( .A(A[6]), .B(n978), .Z(n815) );
  XOR2_X2 U726 ( .A(A[4]), .B(n976), .Z(n816) );
  XOR2_X2 U729 ( .A(A[2]), .B(n974), .Z(n817) );
  XOR2_X2 U732 ( .A(A[0]), .B(n972), .Z(n818) );
  AOI21_X2 U737 ( .B1(n91), .B2(n958), .A(n88), .ZN(n86) );
  XOR2_X2 U738 ( .A(n251), .B(n244), .Z(n937) );
  XOR2_X2 U739 ( .A(n83), .B(n937), .Z(MAC[25]) );
  NAND2_X2 U740 ( .A1(n251), .A2(n83), .ZN(n938) );
  NAND2_X2 U741 ( .A1(n244), .A2(n83), .ZN(n939) );
  NAND2_X2 U742 ( .A1(n244), .A2(n251), .ZN(n940) );
  NAND3_X2 U743 ( .A1(n940), .A2(n939), .A3(n938), .ZN(n82) );
  XOR2_X2 U744 ( .A(n390), .B(n392), .Z(n941) );
  XOR2_X2 U745 ( .A(n388), .B(n941), .Z(n384) );
  NAND2_X2 U746 ( .A1(n390), .A2(n388), .ZN(n942) );
  NAND2_X2 U747 ( .A1(n392), .A2(n388), .ZN(n943) );
  NAND2_X2 U748 ( .A1(n392), .A2(n390), .ZN(n944) );
  NAND3_X2 U749 ( .A1(n944), .A2(n943), .A3(n942), .ZN(n383) );
  AOI21_X2 U750 ( .B1(n127), .B2(n119), .A(n120), .ZN(n118) );
  XNOR2_X1 U751 ( .A(n115), .B(n59), .ZN(MAC[17]) );
  XOR2_X1 U752 ( .A(n52), .B(n86), .Z(MAC[24]) );
  XOR2_X1 U753 ( .A(n60), .B(n118), .Z(MAC[16]) );
  XNOR2_X1 U754 ( .A(n978), .B(B[8]), .ZN(n734) );
  XNOR2_X1 U755 ( .A(n978), .B(B[5]), .ZN(n737) );
  INV_X1 U756 ( .A(A[13]), .ZN(n983) );
  XOR2_X2 U757 ( .A(n972), .B(A[2]), .Z(n945) );
  XOR2_X2 U758 ( .A(n974), .B(A[4]), .Z(n946) );
  XOR2_X2 U759 ( .A(n976), .B(A[6]), .Z(n947) );
  XOR2_X2 U760 ( .A(n980), .B(A[10]), .Z(n948) );
  XOR2_X2 U761 ( .A(A[13]), .B(A[14]), .Z(n949) );
  XOR2_X2 U762 ( .A(n982), .B(A[12]), .Z(n950) );
  OR2_X4 U763 ( .A1(n658), .A2(C[0]), .ZN(n951) );
  AND2_X4 U764 ( .A1(n951), .A2(n194), .ZN(MAC[0]) );
  XNOR2_X2 U765 ( .A(n51), .B(n77), .ZN(n953) );
  INV_X4 U766 ( .A(n953), .ZN(MAC[31]) );
  XNOR2_X1 U767 ( .A(A[15]), .B(B[3]), .ZN(n671) );
  XNOR2_X1 U768 ( .A(n976), .B(B[3]), .ZN(n756) );
  XNOR2_X1 U769 ( .A(n972), .B(B[3]), .ZN(n790) );
  XNOR2_X1 U770 ( .A(n974), .B(B[3]), .ZN(n773) );
  XNOR2_X1 U771 ( .A(A[13]), .B(B[3]), .ZN(n688) );
  XNOR2_X1 U772 ( .A(n978), .B(B[3]), .ZN(n739) );
  XNOR2_X1 U773 ( .A(n982), .B(B[3]), .ZN(n705) );
  XNOR2_X1 U774 ( .A(n980), .B(B[3]), .ZN(n722) );
  AOI21_X2 U775 ( .B1(n115), .B2(n955), .A(n112), .ZN(n110) );
  AOI21_X2 U776 ( .B1(n107), .B2(n956), .A(n104), .ZN(n102) );
  AOI21_X2 U777 ( .B1(n99), .B2(n957), .A(n96), .ZN(n94) );
  NAND2_X2 U778 ( .A1(n816), .A2(n965), .ZN(n18) );
  NAND2_X2 U779 ( .A1(n812), .A2(n969), .ZN(n42) );
  INV_X4 U780 ( .A(n947), .ZN(n966) );
  INV_X4 U781 ( .A(n949), .ZN(n970) );
  INV_X4 U782 ( .A(n973), .ZN(n974) );
  INV_X4 U783 ( .A(n981), .ZN(n982) );
  INV_X2 U784 ( .A(n145), .ZN(n144) );
  NOR2_X1 U785 ( .A1(n121), .A2(n124), .ZN(n119) );
  INV_X1 U786 ( .A(n148), .ZN(n209) );
  INV_X2 U787 ( .A(n143), .ZN(n141) );
  NOR2_X1 U788 ( .A1(n420), .A2(n431), .ZN(n142) );
  NAND2_X1 U789 ( .A1(n432), .A2(n441), .ZN(n149) );
  OAI22_X1 U790 ( .A1(n778), .A2(n6), .B1(n778), .B2(n834), .ZN(n512) );
  OAI22_X1 U791 ( .A1(n42), .A2(n682), .B1(n969), .B2(n681), .ZN(n546) );
  OAI22_X1 U792 ( .A1(n48), .A2(n665), .B1(n970), .B2(n664), .ZN(n529) );
  OAI21_X1 U793 ( .B1(n126), .B2(n124), .A(n125), .ZN(n123) );
  NAND2_X1 U794 ( .A1(n204), .A2(n122), .ZN(n61) );
  OAI22_X1 U795 ( .A1(n676), .A2(n42), .B1(n676), .B2(n969), .ZN(n494) );
  AOI21_X1 U796 ( .B1(n144), .B2(n135), .A(n136), .ZN(n134) );
  NAND2_X1 U797 ( .A1(n954), .A2(n133), .ZN(n63) );
  NAND2_X1 U798 ( .A1(n208), .A2(n143), .ZN(n65) );
  OAI22_X1 U799 ( .A1(n6), .A2(n791), .B1(n790), .B2(n834), .ZN(n655) );
  OAI21_X2 U800 ( .B1(n121), .B2(n125), .A(n122), .ZN(n120) );
  AOI21_X2 U801 ( .B1(n146), .B2(n154), .A(n147), .ZN(n145) );
  NOR2_X2 U802 ( .A1(n148), .A2(n151), .ZN(n146) );
  OAI21_X2 U803 ( .B1(n148), .B2(n152), .A(n149), .ZN(n147) );
  OAI21_X2 U804 ( .B1(n145), .B2(n128), .A(n129), .ZN(n127) );
  AOI21_X2 U805 ( .B1(n954), .B2(n136), .A(n131), .ZN(n129) );
  OAI21_X2 U806 ( .B1(n118), .B2(n116), .A(n117), .ZN(n115) );
  OAI21_X2 U807 ( .B1(n110), .B2(n108), .A(n109), .ZN(n107) );
  OAI21_X2 U808 ( .B1(n102), .B2(n100), .A(n101), .ZN(n99) );
  OAI21_X2 U809 ( .B1(n94), .B2(n92), .A(n93), .ZN(n91) );
  OAI21_X2 U810 ( .B1(n137), .B2(n143), .A(n138), .ZN(n136) );
  OAI21_X2 U811 ( .B1(n157), .B2(n155), .A(n156), .ZN(n154) );
  NOR2_X2 U812 ( .A1(n137), .A2(n142), .ZN(n135) );
  AOI21_X2 U813 ( .B1(n162), .B2(n962), .A(n159), .ZN(n157) );
  AOI21_X2 U814 ( .B1(n959), .B2(n180), .A(n177), .ZN(n175) );
  OAI21_X2 U815 ( .B1(n163), .B2(n175), .A(n164), .ZN(n162) );
  AOI21_X2 U816 ( .B1(n960), .B2(n171), .A(n166), .ZN(n164) );
  NOR2_X2 U817 ( .A1(n408), .A2(n419), .ZN(n137) );
  NOR2_X2 U818 ( .A1(n364), .A2(n379), .ZN(n121) );
  NOR2_X2 U819 ( .A1(n432), .A2(n441), .ZN(n148) );
  NOR2_X2 U820 ( .A1(n380), .A2(n393), .ZN(n124) );
  NOR2_X2 U821 ( .A1(n442), .A2(n451), .ZN(n151) );
  NOR2_X2 U822 ( .A1(n348), .A2(n363), .ZN(n116) );
  NOR2_X2 U823 ( .A1(n318), .A2(n331), .ZN(n108) );
  NOR2_X2 U824 ( .A1(n452), .A2(n459), .ZN(n155) );
  OR2_X1 U825 ( .A1(n394), .A2(n407), .ZN(n954) );
  OR2_X1 U826 ( .A1(n332), .A2(n347), .ZN(n955) );
  OR2_X1 U827 ( .A1(n304), .A2(n317), .ZN(n956) );
  NOR2_X2 U828 ( .A1(n292), .A2(n303), .ZN(n100) );
  NOR2_X2 U829 ( .A1(n270), .A2(n279), .ZN(n92) );
  OR2_X1 U830 ( .A1(n280), .A2(n291), .ZN(n957) );
  OR2_X1 U831 ( .A1(n260), .A2(n269), .ZN(n958) );
  NOR2_X2 U832 ( .A1(n252), .A2(n259), .ZN(n84) );
  OAI21_X2 U833 ( .B1(n181), .B2(n183), .A(n182), .ZN(n180) );
  OAI21_X2 U834 ( .B1(n86), .B2(n84), .A(n85), .ZN(n83) );
  OR2_X1 U835 ( .A1(n480), .A2(n483), .ZN(n959) );
  OR2_X1 U836 ( .A1(n468), .A2(n473), .ZN(n960) );
  OR2_X1 U837 ( .A1(n474), .A2(n479), .ZN(n961) );
  OR2_X1 U838 ( .A1(n460), .A2(n467), .ZN(n962) );
  AOI21_X2 U839 ( .B1(n963), .B2(n192), .A(n189), .ZN(n187) );
  OAI21_X2 U840 ( .B1(n187), .B2(n185), .A(n186), .ZN(n184) );
  INV_X4 U841 ( .A(n512), .ZN(n642) );
  INV_X4 U842 ( .A(n509), .ZN(n625) );
  NOR2_X2 U843 ( .A1(n484), .A2(n486), .ZN(n181) );
  INV_X4 U844 ( .A(n506), .ZN(n608) );
  NOR2_X2 U845 ( .A1(n488), .A2(n489), .ZN(n185) );
  OR2_X1 U846 ( .A1(n490), .A2(n522), .ZN(n963) );
  INV_X4 U847 ( .A(n503), .ZN(n591) );
  INV_X4 U848 ( .A(n500), .ZN(n574) );
  INV_X4 U849 ( .A(n497), .ZN(n557) );
  INV_X4 U850 ( .A(n494), .ZN(n540) );
  AOI21_X2 U851 ( .B1(n144), .B2(n208), .A(n141), .ZN(n139) );
  AOI21_X2 U852 ( .B1(n174), .B2(n961), .A(n171), .ZN(n169) );
  OAI21_X2 U853 ( .B1(n153), .B2(n151), .A(n152), .ZN(n150) );
  XNOR2_X2 U854 ( .A(C[31]), .B(n221), .ZN(n51) );
  NAND2_X2 U855 ( .A1(n815), .A2(n966), .ZN(n24) );
  NAND2_X2 U856 ( .A1(n814), .A2(n28), .ZN(n30) );
  NAND2_X2 U857 ( .A1(n813), .A2(n968), .ZN(n36) );
  NAND2_X2 U858 ( .A1(n811), .A2(n970), .ZN(n48) );
  NAND2_X2 U859 ( .A1(n817), .A2(n964), .ZN(n12) );
  NAND2_X2 U860 ( .A1(n818), .A2(n834), .ZN(n6) );
  INV_X4 U861 ( .A(A[0]), .ZN(n834) );
  INV_X4 U862 ( .A(A[15]), .ZN(n984) );
  INV_X4 U863 ( .A(n979), .ZN(n980) );
  INV_X4 U864 ( .A(A[9]), .ZN(n979) );
  INV_X4 U865 ( .A(n977), .ZN(n978) );
  INV_X4 U866 ( .A(A[7]), .ZN(n977) );
  INV_X4 U867 ( .A(n971), .ZN(n972) );
  INV_X4 U868 ( .A(A[1]), .ZN(n971) );
  INV_X4 U869 ( .A(n975), .ZN(n976) );
  INV_X4 U870 ( .A(A[5]), .ZN(n975) );
  INV_X4 U871 ( .A(A[11]), .ZN(n981) );
  INV_X4 U872 ( .A(A[3]), .ZN(n973) );
  INV_X4 U873 ( .A(n948), .ZN(n968) );
  INV_X4 U874 ( .A(n945), .ZN(n964) );
  INV_X4 U875 ( .A(n28), .ZN(n967) );
  INV_X4 U876 ( .A(n950), .ZN(n969) );
  INV_X4 U877 ( .A(n946), .ZN(n965) );
  INV_X4 U878 ( .A(n491), .ZN(n523) );
  INV_X4 U879 ( .A(n98), .ZN(n96) );
  INV_X4 U880 ( .A(n90), .ZN(n88) );
  OAI22_X2 U881 ( .A1(n761), .A2(n12), .B1(n761), .B2(n964), .ZN(n509) );
  OAI22_X2 U882 ( .A1(n744), .A2(n18), .B1(n744), .B2(n965), .ZN(n506) );
  OAI22_X2 U883 ( .A1(n727), .A2(n24), .B1(n727), .B2(n966), .ZN(n503) );
  OAI22_X2 U884 ( .A1(n710), .A2(n30), .B1(n710), .B2(n28), .ZN(n500) );
  OAI22_X2 U885 ( .A1(n693), .A2(n36), .B1(n693), .B2(n968), .ZN(n497) );
  OAI22_X2 U886 ( .A1(n659), .A2(n48), .B1(n659), .B2(n970), .ZN(n491) );
  INV_X4 U887 ( .A(C[17]), .ZN(n346) );
  INV_X4 U888 ( .A(C[19]), .ZN(n316) );
  INV_X4 U889 ( .A(C[21]), .ZN(n290) );
  INV_X4 U890 ( .A(C[23]), .ZN(n268) );
  INV_X4 U891 ( .A(C[25]), .ZN(n250) );
  INV_X4 U892 ( .A(C[27]), .ZN(n236) );
  INV_X4 U893 ( .A(C[29]), .ZN(n226) );
  INV_X4 U894 ( .A(n185), .ZN(n217) );
  INV_X4 U895 ( .A(n181), .ZN(n216) );
  INV_X4 U896 ( .A(n155), .ZN(n211) );
  INV_X4 U897 ( .A(n151), .ZN(n210) );
  INV_X4 U898 ( .A(n137), .ZN(n207) );
  INV_X4 U899 ( .A(n124), .ZN(n205) );
  INV_X4 U900 ( .A(n121), .ZN(n204) );
  INV_X4 U901 ( .A(n116), .ZN(n203) );
  INV_X4 U902 ( .A(n108), .ZN(n201) );
  INV_X4 U903 ( .A(n100), .ZN(n199) );
  INV_X4 U904 ( .A(n92), .ZN(n197) );
  INV_X4 U905 ( .A(n84), .ZN(n195) );
  INV_X4 U906 ( .A(n194), .ZN(n192) );
  INV_X4 U907 ( .A(n191), .ZN(n189) );
  INV_X4 U908 ( .A(n184), .ZN(n183) );
  INV_X4 U909 ( .A(n179), .ZN(n177) );
  INV_X4 U910 ( .A(n175), .ZN(n174) );
  INV_X4 U911 ( .A(n173), .ZN(n171) );
  INV_X4 U912 ( .A(n168), .ZN(n166) );
  INV_X4 U913 ( .A(n161), .ZN(n159) );
  INV_X4 U914 ( .A(n154), .ZN(n153) );
  INV_X4 U915 ( .A(n142), .ZN(n208) );
  INV_X4 U916 ( .A(n133), .ZN(n131) );
  INV_X4 U917 ( .A(n127), .ZN(n126) );
  INV_X4 U918 ( .A(n114), .ZN(n112) );
  INV_X4 U919 ( .A(n106), .ZN(n104) );
endmodule


module macopertion_2 ( in_a_mac, in_b_mac, bitselect1, clk, min );
  input [15:0] in_a_mac;
  input [15:0] in_b_mac;
  input [3:0] bitselect1;
  output [15:0] min;
  input clk;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18,
         N19, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49,
         N50, N51, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197;
  wire   [31:0] in_c_mac;
  wire   [31:0] out_mac;
  assign min[15] = 1'b0;

  macopertion_2_DW02_mac_1 U1 ( .A(in_a_mac), .B({in_b_mac[15:1], n179}), .C(
        in_c_mac), .TC(1'b1), .MAC(out_mac) );
  DFF_X1 in_c_mac_reg_0_ ( .D(N4), .CK(clk), .Q(in_c_mac[0]) );
  DFF_X1 in_c_mac_reg_1_ ( .D(N5), .CK(clk), .Q(in_c_mac[1]) );
  DFF_X1 in_c_mac_reg_2_ ( .D(N6), .CK(clk), .Q(in_c_mac[2]) );
  DFF_X1 in_c_mac_reg_3_ ( .D(N7), .CK(clk), .Q(in_c_mac[3]) );
  DFF_X1 in_c_mac_reg_4_ ( .D(N8), .CK(clk), .Q(in_c_mac[4]) );
  DFF_X1 in_c_mac_reg_5_ ( .D(N9), .CK(clk), .Q(in_c_mac[5]) );
  DFF_X1 in_c_mac_reg_6_ ( .D(N10), .CK(clk), .Q(in_c_mac[6]) );
  DFF_X1 in_c_mac_reg_7_ ( .D(N11), .CK(clk), .Q(in_c_mac[7]) );
  DFF_X1 in_c_mac_reg_8_ ( .D(N12), .CK(clk), .Q(in_c_mac[8]) );
  DFF_X1 in_c_mac_reg_9_ ( .D(N13), .CK(clk), .Q(in_c_mac[9]) );
  DFF_X1 in_c_mac_reg_10_ ( .D(N14), .CK(clk), .Q(in_c_mac[10]) );
  DFF_X1 in_c_mac_reg_11_ ( .D(N15), .CK(clk), .Q(in_c_mac[11]) );
  DFF_X1 in_c_mac_reg_12_ ( .D(N16), .CK(clk), .Q(in_c_mac[12]) );
  DFF_X1 in_c_mac_reg_13_ ( .D(N17), .CK(clk), .Q(in_c_mac[13]) );
  DFF_X1 in_c_mac_reg_14_ ( .D(N18), .CK(clk), .Q(in_c_mac[14]) );
  DFF_X1 in_c_mac_reg_15_ ( .D(N19), .CK(clk), .Q(in_c_mac[15]) );
  SDFF_X1 in_c_mac_reg_16_ ( .D(out_mac[16]), .SI(1'b0), .SE(n197), .CK(clk), 
        .Q(in_c_mac[16]) );
  SDFF_X1 in_c_mac_reg_17_ ( .D(out_mac[17]), .SI(1'b0), .SE(n197), .CK(clk), 
        .Q(in_c_mac[17]) );
  SDFF_X1 in_c_mac_reg_18_ ( .D(out_mac[18]), .SI(1'b0), .SE(n197), .CK(clk), 
        .Q(in_c_mac[18]) );
  SDFF_X1 in_c_mac_reg_19_ ( .D(out_mac[19]), .SI(1'b0), .SE(n197), .CK(clk), 
        .Q(in_c_mac[19]) );
  SDFF_X1 in_c_mac_reg_20_ ( .D(out_mac[20]), .SI(1'b0), .SE(n197), .CK(clk), 
        .Q(in_c_mac[20]) );
  SDFF_X1 in_c_mac_reg_21_ ( .D(out_mac[21]), .SI(1'b0), .SE(n197), .CK(clk), 
        .Q(in_c_mac[21]) );
  SDFF_X1 in_c_mac_reg_22_ ( .D(out_mac[22]), .SI(1'b0), .SE(n197), .CK(clk), 
        .Q(in_c_mac[22]) );
  SDFF_X1 in_c_mac_reg_23_ ( .D(out_mac[23]), .SI(1'b0), .SE(n197), .CK(clk), 
        .Q(in_c_mac[23]) );
  SDFF_X1 in_c_mac_reg_24_ ( .D(out_mac[24]), .SI(1'b0), .SE(n197), .CK(clk), 
        .Q(in_c_mac[24]) );
  SDFF_X1 in_c_mac_reg_25_ ( .D(out_mac[25]), .SI(1'b0), .SE(n197), .CK(clk), 
        .Q(in_c_mac[25]) );
  SDFF_X1 in_c_mac_reg_26_ ( .D(out_mac[26]), .SI(1'b0), .SE(n197), .CK(clk), 
        .Q(in_c_mac[26]) );
  SDFF_X1 in_c_mac_reg_27_ ( .D(out_mac[27]), .SI(1'b0), .SE(n197), .CK(clk), 
        .Q(in_c_mac[27]) );
  SDFF_X1 in_c_mac_reg_28_ ( .D(out_mac[28]), .SI(1'b0), .SE(n197), .CK(clk), 
        .Q(in_c_mac[28]) );
  SDFF_X1 in_c_mac_reg_29_ ( .D(out_mac[29]), .SI(1'b0), .SE(n197), .CK(clk), 
        .Q(in_c_mac[29]) );
  SDFF_X1 in_c_mac_reg_30_ ( .D(out_mac[30]), .SI(1'b0), .SE(n197), .CK(clk), 
        .Q(in_c_mac[30]) );
  DFF_X1 min_reg_14_ ( .D(N51), .CK(clk), .Q(min[14]) );
  DFF_X1 min_reg_13_ ( .D(N50), .CK(clk), .Q(min[13]) );
  DFF_X1 min_reg_12_ ( .D(N49), .CK(clk), .Q(min[12]) );
  DFF_X1 min_reg_11_ ( .D(N48), .CK(clk), .Q(min[11]) );
  DFF_X1 min_reg_10_ ( .D(N47), .CK(clk), .Q(min[10]) );
  DFF_X1 min_reg_9_ ( .D(N46), .CK(clk), .Q(min[9]) );
  DFF_X1 min_reg_8_ ( .D(N45), .CK(clk), .Q(min[8]) );
  DFF_X1 min_reg_7_ ( .D(N44), .CK(clk), .Q(min[7]) );
  DFF_X1 min_reg_6_ ( .D(N43), .CK(clk), .Q(min[6]) );
  DFF_X1 min_reg_5_ ( .D(N42), .CK(clk), .Q(min[5]) );
  DFF_X1 min_reg_4_ ( .D(N41), .CK(clk), .Q(min[4]) );
  DFF_X1 min_reg_3_ ( .D(N40), .CK(clk), .Q(min[3]) );
  DFF_X1 min_reg_2_ ( .D(N39), .CK(clk), .Q(min[2]) );
  DFF_X1 min_reg_1_ ( .D(N38), .CK(clk), .Q(min[1]) );
  DFF_X1 min_reg_0_ ( .D(N37), .CK(clk), .Q(min[0]) );
  SDFF_X2 in_c_mac_reg_31_ ( .D(out_mac[31]), .SI(1'b0), .SE(n197), .CK(clk), 
        .Q(in_c_mac[31]) );
  INV_X4 U23 ( .A(n180), .ZN(n179) );
  INV_X1 U24 ( .A(in_b_mac[0]), .ZN(n180) );
  INV_X4 U25 ( .A(n181), .ZN(n197) );
  OR4_X4 U26 ( .A1(bitselect1[1]), .A2(bitselect1[0]), .A3(bitselect1[3]), 
        .A4(bitselect1[2]), .ZN(n181) );
  AND2_X1 U27 ( .A1(out_mac[15]), .A2(n181), .ZN(N19) );
  AND2_X1 U28 ( .A1(out_mac[14]), .A2(n181), .ZN(N18) );
  AND2_X1 U29 ( .A1(out_mac[13]), .A2(n181), .ZN(N17) );
  AND2_X1 U30 ( .A1(out_mac[12]), .A2(n181), .ZN(N16) );
  AND2_X1 U31 ( .A1(out_mac[11]), .A2(n181), .ZN(N15) );
  AND2_X1 U32 ( .A1(out_mac[10]), .A2(n181), .ZN(N14) );
  AND2_X1 U33 ( .A1(out_mac[9]), .A2(n181), .ZN(N13) );
  AND2_X1 U34 ( .A1(out_mac[8]), .A2(n181), .ZN(N12) );
  AND2_X1 U35 ( .A1(out_mac[7]), .A2(n181), .ZN(N11) );
  AND2_X1 U36 ( .A1(out_mac[6]), .A2(n181), .ZN(N10) );
  AND2_X1 U37 ( .A1(out_mac[5]), .A2(n181), .ZN(N9) );
  AND2_X1 U38 ( .A1(out_mac[4]), .A2(n181), .ZN(N8) );
  AND2_X1 U39 ( .A1(out_mac[3]), .A2(n181), .ZN(N7) );
  AND2_X1 U40 ( .A1(out_mac[2]), .A2(n181), .ZN(N6) );
  AND2_X1 U41 ( .A1(out_mac[1]), .A2(n181), .ZN(N5) );
  AND2_X1 U42 ( .A1(out_mac[0]), .A2(n181), .ZN(N4) );
  INV_X4 U43 ( .A(out_mac[16]), .ZN(n182) );
  NOR2_X2 U44 ( .A1(out_mac[31]), .A2(n182), .ZN(N37) );
  INV_X4 U45 ( .A(out_mac[17]), .ZN(n183) );
  NOR2_X2 U46 ( .A1(out_mac[31]), .A2(n183), .ZN(N38) );
  INV_X4 U47 ( .A(out_mac[18]), .ZN(n184) );
  NOR2_X2 U48 ( .A1(out_mac[31]), .A2(n184), .ZN(N39) );
  INV_X4 U49 ( .A(out_mac[19]), .ZN(n185) );
  NOR2_X2 U50 ( .A1(out_mac[31]), .A2(n185), .ZN(N40) );
  INV_X4 U51 ( .A(out_mac[20]), .ZN(n186) );
  NOR2_X2 U52 ( .A1(out_mac[31]), .A2(n186), .ZN(N41) );
  INV_X4 U53 ( .A(out_mac[21]), .ZN(n187) );
  NOR2_X2 U54 ( .A1(out_mac[31]), .A2(n187), .ZN(N42) );
  INV_X4 U55 ( .A(out_mac[22]), .ZN(n188) );
  NOR2_X2 U56 ( .A1(out_mac[31]), .A2(n188), .ZN(N43) );
  INV_X4 U57 ( .A(out_mac[23]), .ZN(n189) );
  NOR2_X2 U58 ( .A1(out_mac[31]), .A2(n189), .ZN(N44) );
  INV_X4 U59 ( .A(out_mac[24]), .ZN(n190) );
  NOR2_X2 U60 ( .A1(out_mac[31]), .A2(n190), .ZN(N45) );
  INV_X4 U61 ( .A(out_mac[25]), .ZN(n191) );
  NOR2_X2 U62 ( .A1(out_mac[31]), .A2(n191), .ZN(N46) );
  INV_X4 U63 ( .A(out_mac[26]), .ZN(n192) );
  NOR2_X2 U64 ( .A1(out_mac[31]), .A2(n192), .ZN(N47) );
  INV_X4 U65 ( .A(out_mac[27]), .ZN(n193) );
  NOR2_X2 U66 ( .A1(out_mac[31]), .A2(n193), .ZN(N48) );
  INV_X4 U67 ( .A(out_mac[28]), .ZN(n194) );
  NOR2_X2 U68 ( .A1(out_mac[31]), .A2(n194), .ZN(N49) );
  INV_X4 U69 ( .A(out_mac[29]), .ZN(n195) );
  NOR2_X2 U70 ( .A1(out_mac[31]), .A2(n195), .ZN(N50) );
  INV_X4 U71 ( .A(out_mac[30]), .ZN(n196) );
  NOR2_X2 U72 ( .A1(out_mac[31]), .A2(n196), .ZN(N51) );
endmodule


module macopertion_0 ( in_a_mac, in_b_mac, bitselect1, clk, min );
  input [15:0] in_a_mac;
  input [15:0] in_b_mac;
  input [3:0] bitselect1;
  output [15:0] min;
  input clk;
  wire   U6_Z_0, U6_Z_1, U6_Z_2, U6_Z_3, U6_Z_4, U6_Z_5, U6_Z_6, U6_Z_7,
         U6_Z_8, U6_Z_9, U6_Z_10, U6_Z_11, U6_Z_12, U6_Z_13, U6_Z_14, U6_Z_15,
         U6_Z_16, U6_Z_17, U6_Z_18, U6_Z_19, U6_Z_20, U6_Z_21, U6_Z_22,
         U6_Z_23, U6_Z_24, U6_Z_25, U6_Z_26, U6_Z_27, U6_Z_28, U6_Z_29,
         U6_Z_30, U5_Z_0, U5_Z_1, U5_Z_2, U5_Z_3, U5_Z_4, U5_Z_5, U5_Z_6,
         U5_Z_7, U5_Z_8, U5_Z_9, U5_Z_10, U5_Z_11, U5_Z_12, U5_Z_13, U5_Z_14,
         U1_C_31_, U1_C_30_, U1_C_28_, U1_C_26_, U1_C_24_, U1_C_22_, U1_C_20_,
         U1_C_18_, U1_C_16_, U1_C_15_, U1_C_14_, U1_C_13_, U1_C_12_, U1_C_11_,
         U1_C_10_, U1_C_9_, U1_C_8_, U1_C_7_, U1_C_6_, U1_C_5_, U1_C_4_,
         U1_C_3_, U1_C_2_, U1_C_1_, U1_C_0_, U1_C_17_, U1_C_21_, U1_C_23_,
         U1_C_25_, U1_C_27_, n4, n12, n18, n29, n41, n52, n65, n208, n209,
         n212, n217, n242, n243, n244, n245, n247, n248, n249, n250, n255,
         n256, n257, n258, n259, n264, n269, n274, n279, n283, n360, n361,
         n362, n366, n367, n368, n559, n574, n590, n595, n596, n613, n614,
         n616, n621, n623, n624, n635, n640, n642, n644, n646, n647, n653,
         n656, n657, n660, n661, n664, n665, n672, n673, n674, n675, n676,
         n684, n686, n688, n691, n692, n696, n698, n700, n701, n706, n707,
         n708, n709, n710, n714, n720, n721, n722, n724, n725, n726, n729,
         n731, n732, n733, n735, n739, n740, n746, n747, n750, n751, n754,
         n756, n757, n760, n762, n764, n765, n766, n769, n770, n774, n775,
         n776, n777, n779, n783, n789, n791, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n820, n821, n822,
         n823, n825, n826, n829, n830, n833, n835, n836, n837, n838, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n852, n854,
         n860, n861, n862, n864, n868, n869, n870, n871, n872, n873, n874,
         n876, n878, n879, n881, n883, n884, n885, n886, n887, n888, n889,
         n890, n892, n893, n895, n896, n897, n898, n899, n900, n903, n905,
         n907, n908, n909, n910, n911, n912, n913, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n935, n937, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n954, n956, n957, n958, n959, n960, n962, n963, n964,
         n965, n966, n967, n970, n971, n972, n973, n975, n976, n978, n979,
         n980, n982, n983, n984, n986, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1003, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1016, n1018, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1041, n1042,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1091, n1092, n1093, n1094, n1095, n1096,
         n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1119, n1120, n1121, n1122, n1123, n1124, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n210, n211, n213, n214, n215, n216, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n246, n251, n252, n253, n254, n260, n261, n262, n263, n265, n266,
         n267, n268, n270, n271, n272, n273, n275, n276, n277, n278, n280,
         n281, n282, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n363, n364, n365, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n591, n592, n593, n594, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n615, n617, n618, n619, n620, n622, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n636, n637, n638, n639, n641,
         n643, n645, n648, n649, n650, n651, n652, n654, n655, n658, n659,
         n662, n663, n666, n667, n668, n669, n670, n671, n677, n678, n679,
         n680, n681, n682, n683, n685, n687, n689, n690, n693, n694, n695,
         n697, n699, n702, n703, n704, n705, n711, n712, n713, n715, n716,
         n717, n718, n719, n723, n727, n728, n730, n734, n736, n737, n738,
         n741, n742, n743, n744, n745, n748, n749, n752, n753, n755, n758,
         n759, n761, n763, n767, n768, n771, n772, n773, n778, n780, n781,
         n782, n784, n785, n786, n787, n788, n790, n792, n807, n818, n819,
         n824, n827, n828, n831, n832, n834, n839, n850, n851, n853, n855,
         n856, n857, n858, n859, n863, n865, n866, n867, n875, n877, n880,
         n882, n891, n894, n901, n902, n904, n906, n914, n915, n916, n917,
         n933, n934, n936, n938, n950, n951, n952, n953, n955, n961, n968,
         n969, n974, n977, n981, n985, n987, n1002, n1004, n1005, n1014, n1015,
         n1017, n1019, n1040, n1043, n1044, n1073, n1090, n1106, n1118, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
         n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
         n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
         n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
         n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
         n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
         n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
         n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554;
  assign min[15] = 1'b0;

  NOR2_X2 U6 ( .A1(n208), .A2(n209), .ZN(U6_Z_9) );
  NOR2_X2 U9 ( .A1(n208), .A2(n212), .ZN(U6_Z_8) );
  NOR2_X2 U12 ( .A1(n208), .A2(n217), .ZN(U6_Z_7) );
  NOR2_X2 U29 ( .A1(n208), .A2(n242), .ZN(U6_Z_28) );
  NOR2_X2 U30 ( .A1(n208), .A2(n243), .ZN(U6_Z_27) );
  NOR2_X2 U31 ( .A1(n208), .A2(n244), .ZN(U6_Z_26) );
  NOR2_X2 U32 ( .A1(n208), .A2(n245), .ZN(U6_Z_25) );
  NOR2_X2 U35 ( .A1(n208), .A2(n248), .ZN(U6_Z_22) );
  NOR2_X2 U36 ( .A1(n208), .A2(n249), .ZN(U6_Z_21) );
  NOR2_X2 U37 ( .A1(n208), .A2(n250), .ZN(U6_Z_20) );
  NOR2_X2 U41 ( .A1(n208), .A2(n255), .ZN(U6_Z_19) );
  NOR2_X2 U42 ( .A1(n208), .A2(n256), .ZN(U6_Z_18) );
  NOR2_X2 U43 ( .A1(n208), .A2(n257), .ZN(U6_Z_17) );
  NOR2_X2 U44 ( .A1(n208), .A2(n258), .ZN(U6_Z_16) );
  NOR2_X2 U45 ( .A1(n208), .A2(n259), .ZN(U6_Z_15) );
  NOR2_X2 U48 ( .A1(n208), .A2(n264), .ZN(U6_Z_14) );
  NOR2_X2 U51 ( .A1(n208), .A2(n269), .ZN(U6_Z_13) );
  NOR2_X2 U54 ( .A1(n208), .A2(n274), .ZN(U6_Z_12) );
  NOR2_X2 U57 ( .A1(n208), .A2(n279), .ZN(U6_Z_11) );
  NOR2_X2 U60 ( .A1(n208), .A2(n283), .ZN(U6_Z_10) );
  XOR2_X2 U132 ( .A(in_b_mac[15]), .B(n1554), .Z(n362) );
  XNOR2_X2 U329 ( .A(in_b_mac[6]), .B(n434), .ZN(n574) );
  XNOR2_X2 U350 ( .A(in_b_mac[7]), .B(n434), .ZN(n590) );
  XOR2_X2 U354 ( .A(in_b_mac[1]), .B(n1551), .Z(n595) );
  XNOR2_X2 U393 ( .A(in_b_mac[8]), .B(n434), .ZN(n614) );
  XOR2_X2 U401 ( .A(in_b_mac[2]), .B(n1551), .Z(n616) );
  OAI22_X2 U421 ( .A1(n440), .A2(n691), .B1(n640), .B2(n642), .ZN(n635) );
  XNOR2_X2 U422 ( .A(in_b_mac[1]), .B(n436), .ZN(n640) );
  XNOR2_X2 U440 ( .A(n708), .B(n1547), .ZN(n674) );
  XOR2_X2 U441 ( .A(n709), .B(n710), .Z(n708) );
  OAI22_X2 U453 ( .A1(n440), .A2(n722), .B1(n691), .B2(n280), .ZN(n656) );
  XNOR2_X2 U454 ( .A(in_b_mac[2]), .B(n436), .ZN(n691) );
  OAI22_X2 U457 ( .A1(n438), .A2(n724), .B1(n725), .B2(n721), .ZN(n653) );
  XOR2_X2 U458 ( .A(n1552), .B(n443), .Z(n725) );
  XOR2_X2 U460 ( .A(in_b_mac[4]), .B(n1551), .Z(n692) );
  OAI22_X2 U486 ( .A1(n438), .A2(n756), .B1(n724), .B2(n721), .ZN(n686) );
  XOR2_X2 U487 ( .A(in_b_mac[1]), .B(n1552), .Z(n724) );
  XOR2_X2 U495 ( .A(in_b_mac[5]), .B(n1551), .Z(n726) );
  XOR2_X2 U530 ( .A(n795), .B(n796), .Z(n766) );
  XOR2_X2 U531 ( .A(n797), .B(n798), .Z(n796) );
  XOR2_X2 U534 ( .A(n800), .B(n801), .Z(n729) );
  XOR2_X2 U535 ( .A(n802), .B(n803), .Z(n801) );
  XOR2_X2 U536 ( .A(n804), .B(n805), .Z(n732) );
  OAI22_X2 U542 ( .A1(n437), .A2(n812), .B1(n813), .B2(n814), .ZN(n710) );
  XNOR2_X2 U546 ( .A(in_b_mac[4]), .B(n230), .ZN(n757) );
  XOR2_X2 U555 ( .A(in_b_mac[6]), .B(n1551), .Z(n760) );
  OAI22_X2 U556 ( .A1(n438), .A2(n821), .B1(n756), .B2(n721), .ZN(n754) );
  XOR2_X2 U557 ( .A(in_b_mac[2]), .B(n1552), .Z(n756) );
  OAI22_X2 U562 ( .A1(n437), .A2(n825), .B1(n812), .B2(n814), .ZN(n779) );
  XOR2_X2 U563 ( .A(in_b_mac[1]), .B(n1553), .Z(n812) );
  OAI22_X2 U564 ( .A1(n438), .A2(n826), .B1(n821), .B2(n721), .ZN(n777) );
  XOR2_X2 U565 ( .A(n320), .B(n1552), .Z(n821) );
  XNOR2_X2 U571 ( .A(in_b_mac[5]), .B(n230), .ZN(n816) );
  XOR2_X2 U573 ( .A(in_b_mac[7]), .B(n1551), .Z(n820) );
  XOR2_X2 U584 ( .A(n837), .B(n838), .Z(n836) );
  XNOR2_X2 U589 ( .A(n1509), .B(n846), .ZN(n793) );
  XNOR2_X2 U590 ( .A(n847), .B(n848), .ZN(n846) );
  XNOR2_X2 U595 ( .A(n1514), .B(n852), .ZN(n765) );
  XNOR2_X2 U596 ( .A(n423), .B(n854), .ZN(n852) );
  XOR2_X2 U603 ( .A(in_b_mac[8]), .B(n1551), .Z(n830) );
  OAI22_X2 U604 ( .A1(n797), .A2(n798), .B1(n861), .B2(n795), .ZN(n843) );
  OAI22_X2 U612 ( .A1(n438), .A2(n869), .B1(n826), .B2(n721), .ZN(n805) );
  XOR2_X2 U613 ( .A(in_b_mac[4]), .B(n1552), .Z(n826) );
  OAI22_X2 U616 ( .A1(n361), .A2(n871), .B1(n872), .B2(n360), .ZN(n802) );
  XNOR2_X2 U619 ( .A(in_b_mac[6]), .B(n230), .ZN(n829) );
  OAI22_X2 U620 ( .A1(n437), .A2(n874), .B1(n825), .B2(n814), .ZN(n803) );
  XOR2_X2 U621 ( .A(n317), .B(n1553), .Z(n825) );
  XOR2_X2 U627 ( .A(n1502), .B(n883), .Z(n881) );
  XNOR2_X2 U630 ( .A(n885), .B(n886), .ZN(n840) );
  XOR2_X2 U631 ( .A(n887), .B(n888), .Z(n886) );
  OAI22_X2 U636 ( .A1(n361), .A2(n892), .B1(n871), .B2(n360), .ZN(n864) );
  XOR2_X2 U637 ( .A(in_b_mac[1]), .B(n1554), .Z(n871) );
  OAI22_X2 U638 ( .A1(n437), .A2(n893), .B1(n874), .B2(n814), .ZN(n862) );
  XOR2_X2 U639 ( .A(n320), .B(n1553), .Z(n874) );
  XNOR2_X2 U648 ( .A(in_b_mac[7]), .B(n230), .ZN(n873) );
  OAI22_X2 U653 ( .A1(n438), .A2(n905), .B1(n869), .B2(n721), .ZN(n903) );
  XOR2_X2 U654 ( .A(in_b_mac[5]), .B(n1552), .Z(n869) );
  XNOR2_X2 U660 ( .A(n908), .B(n909), .ZN(n791) );
  XOR2_X2 U661 ( .A(n910), .B(n911), .Z(n909) );
  XOR2_X2 U662 ( .A(n1513), .B(n912), .Z(n789) );
  XNOR2_X2 U663 ( .A(n913), .B(n1542), .ZN(n912) );
  XOR2_X2 U669 ( .A(n920), .B(n921), .Z(n919) );
  XOR2_X2 U671 ( .A(n1515), .B(n924), .Z(n923) );
  XOR2_X2 U674 ( .A(n928), .B(n929), .Z(n927) );
  XNOR2_X2 U677 ( .A(n931), .B(n932), .ZN(n838) );
  XOR2_X2 U678 ( .A(U1_C_18_), .B(n65), .Z(n931) );
  XOR2_X2 U681 ( .A(n937), .B(n1544), .Z(n837) );
  OAI22_X2 U687 ( .A1(n361), .A2(n942), .B1(n892), .B2(n360), .ZN(n910) );
  XOR2_X2 U688 ( .A(n317), .B(n1554), .Z(n892) );
  OAI22_X2 U689 ( .A1(n437), .A2(n943), .B1(n893), .B2(n814), .ZN(n908) );
  XOR2_X2 U690 ( .A(in_b_mac[4]), .B(n1553), .Z(n893) );
  OAI22_X2 U694 ( .A1(n438), .A2(n948), .B1(n905), .B2(n721), .ZN(n913) );
  XOR2_X2 U695 ( .A(in_b_mac[6]), .B(n1552), .Z(n905) );
  NOR2_X2 U696 ( .A1(n898), .A2(U1_C_16_), .ZN(n899) );
  XOR2_X2 U698 ( .A(in_b_mac[9]), .B(n1551), .Z(n860) );
  XOR2_X2 U699 ( .A(in_b_mac[10]), .B(n1551), .Z(n945) );
  XNOR2_X2 U701 ( .A(in_b_mac[8]), .B(n230), .ZN(n900) );
  XOR2_X2 U713 ( .A(n960), .B(n1520), .Z(n959) );
  XNOR2_X2 U717 ( .A(n965), .B(n966), .ZN(n963) );
  XNOR2_X2 U722 ( .A(n970), .B(n971), .ZN(n879) );
  XOR2_X2 U723 ( .A(n972), .B(n973), .Z(n971) );
  OAI22_X2 U726 ( .A1(n437), .A2(n975), .B1(n943), .B2(n814), .ZN(n935) );
  XOR2_X2 U727 ( .A(in_b_mac[5]), .B(n1553), .Z(n943) );
  XOR2_X2 U729 ( .A(in_b_mac[11]), .B(n1551), .Z(n944) );
  XNOR2_X2 U737 ( .A(in_b_mac[9]), .B(n230), .ZN(n949) );
  OAI22_X2 U740 ( .A1(n361), .A2(n983), .B1(n942), .B2(n360), .ZN(n939) );
  XOR2_X2 U741 ( .A(n320), .B(n1554), .Z(n942) );
  XOR2_X2 U743 ( .A(in_b_mac[7]), .B(n1552), .Z(n948) );
  OAI22_X2 U749 ( .A1(n437), .A2(n986), .B1(n975), .B2(n814), .ZN(n929) );
  XOR2_X2 U750 ( .A(in_b_mac[6]), .B(n1553), .Z(n975) );
  XOR2_X2 U754 ( .A(n990), .B(n1529), .Z(n989) );
  XOR2_X2 U756 ( .A(n993), .B(n994), .Z(n992) );
  XOR2_X2 U759 ( .A(n997), .B(n998), .Z(n958) );
  XOR2_X2 U760 ( .A(n999), .B(n1000), .Z(n998) );
  OAI22_X2 U761 ( .A1(n920), .A2(n921), .B1(n1001), .B2(n918), .ZN(n996) );
  XOR2_X2 U764 ( .A(n1006), .B(n1007), .Z(n921) );
  XNOR2_X2 U765 ( .A(U1_C_20_), .B(n593), .ZN(n1006) );
  OAI22_X2 U768 ( .A1(n361), .A2(n1009), .B1(n983), .B2(n360), .ZN(n972) );
  XOR2_X2 U769 ( .A(in_b_mac[4]), .B(n1554), .Z(n983) );
  OAI22_X2 U770 ( .A1(n438), .A2(n1010), .B1(n984), .B2(n721), .ZN(n970) );
  XOR2_X2 U771 ( .A(in_b_mac[8]), .B(n1552), .Z(n984) );
  XNOR2_X2 U773 ( .A(in_b_mac[10]), .B(n230), .ZN(n980) );
  OAI22_X2 U776 ( .A1(n361), .A2(n1013), .B1(n1009), .B2(n360), .ZN(n966) );
  XOR2_X2 U777 ( .A(in_b_mac[5]), .B(n1554), .Z(n1009) );
  XOR2_X2 U781 ( .A(in_b_mac[12]), .B(n1551), .Z(n976) );
  OAI22_X2 U784 ( .A1(n437), .A2(n1018), .B1(n986), .B2(n814), .ZN(n965) );
  XOR2_X2 U785 ( .A(in_b_mac[7]), .B(n1553), .Z(n986) );
  XNOR2_X2 U789 ( .A(n1022), .B(n1023), .ZN(n1020) );
  XOR2_X2 U791 ( .A(n1026), .B(n1027), .Z(n1025) );
  XOR2_X2 U794 ( .A(n1029), .B(n1533), .Z(n991) );
  XOR2_X2 U795 ( .A(U1_C_22_), .B(n41), .Z(n1029) );
  XNOR2_X2 U796 ( .A(n1030), .B(n1031), .ZN(n994) );
  XOR2_X2 U797 ( .A(n1032), .B(n1033), .Z(n1030) );
  XNOR2_X2 U800 ( .A(n1035), .B(n1036), .ZN(n954) );
  XOR2_X2 U801 ( .A(n41), .B(n1037), .Z(n1036) );
  XNOR2_X2 U805 ( .A(in_b_mac[11]), .B(n230), .ZN(n1011) );
  XOR2_X2 U809 ( .A(in_b_mac[13]), .B(n1551), .Z(n1016) );
  OAI22_X2 U810 ( .A1(n438), .A2(n1042), .B1(n1010), .B2(n721), .ZN(n1003) );
  XOR2_X2 U811 ( .A(in_b_mac[9]), .B(n1552), .Z(n1010) );
  XOR2_X2 U819 ( .A(n1047), .B(n1048), .Z(n1046) );
  XOR2_X2 U822 ( .A(n1050), .B(n1051), .Z(n1024) );
  XOR2_X2 U823 ( .A(n29), .B(n1052), .Z(n1051) );
  XNOR2_X2 U829 ( .A(in_b_mac[12]), .B(n230), .ZN(n1039) );
  XOR2_X2 U831 ( .A(in_b_mac[14]), .B(n1551), .Z(n1041) );
  OAI22_X2 U834 ( .A1(n437), .A2(n1058), .B1(n1018), .B2(n814), .ZN(n999) );
  XOR2_X2 U835 ( .A(in_b_mac[8]), .B(n1553), .Z(n1018) );
  OAI22_X2 U836 ( .A1(n438), .A2(n1059), .B1(n1042), .B2(n721), .ZN(n997) );
  XOR2_X2 U837 ( .A(in_b_mac[10]), .B(n1552), .Z(n1042) );
  OAI22_X2 U838 ( .A1(n361), .A2(n1060), .B1(n1013), .B2(n360), .ZN(n1000) );
  XOR2_X2 U839 ( .A(in_b_mac[6]), .B(n1554), .Z(n1013) );
  XNOR2_X2 U841 ( .A(in_b_mac[13]), .B(n230), .ZN(n1055) );
  OAI22_X2 U844 ( .A1(n361), .A2(n1064), .B1(n1060), .B2(n360), .ZN(n1033) );
  XOR2_X2 U845 ( .A(in_b_mac[7]), .B(n1554), .Z(n1060) );
  OAI22_X2 U846 ( .A1(n437), .A2(n1065), .B1(n1058), .B2(n814), .ZN(n1031) );
  XOR2_X2 U847 ( .A(in_b_mac[9]), .B(n1553), .Z(n1058) );
  XOR2_X2 U849 ( .A(in_b_mac[15]), .B(n1551), .Z(n1056) );
  OAI22_X2 U855 ( .A1(n361), .A2(n1068), .B1(n1064), .B2(n360), .ZN(n1023) );
  XOR2_X2 U856 ( .A(in_b_mac[8]), .B(n1554), .Z(n1064) );
  OAI22_X2 U859 ( .A1(n438), .A2(n1071), .B1(n1059), .B2(n721), .ZN(n1070) );
  XOR2_X2 U860 ( .A(in_b_mac[11]), .B(n1552), .Z(n1059) );
  OAI22_X2 U861 ( .A1(n437), .A2(n1072), .B1(n1065), .B2(n814), .ZN(n1022) );
  XOR2_X2 U862 ( .A(in_b_mac[10]), .B(n1553), .Z(n1065) );
  XOR2_X2 U866 ( .A(n18), .B(n1076), .Z(n1075) );
  XOR2_X2 U868 ( .A(n1079), .B(n1080), .Z(n1078) );
  XOR2_X2 U871 ( .A(n1082), .B(n1083), .Z(n1045) );
  XOR2_X2 U872 ( .A(U1_C_24_), .B(n29), .Z(n1082) );
  XNOR2_X2 U873 ( .A(n1084), .B(n1539), .ZN(n1048) );
  XOR2_X2 U874 ( .A(n1085), .B(n1086), .Z(n1084) );
  OAI22_X2 U877 ( .A1(n438), .A2(n1088), .B1(n1071), .B2(n721), .ZN(n1050) );
  XOR2_X2 U878 ( .A(in_b_mac[12]), .B(n1552), .Z(n1071) );
  XNOR2_X2 U880 ( .A(in_b_mac[14]), .B(n230), .ZN(n1062) );
  XOR2_X2 U884 ( .A(U1_C_26_), .B(n18), .Z(n1091) );
  XOR2_X2 U886 ( .A(n1095), .B(n1096), .Z(n1093) );
  OAI22_X2 U891 ( .A1(n438), .A2(n1099), .B1(n1088), .B2(n721), .ZN(n1083) );
  XOR2_X2 U892 ( .A(in_b_mac[13]), .B(n1552), .Z(n1088) );
  OAI22_X2 U895 ( .A1(n437), .A2(n1102), .B1(n1072), .B2(n814), .ZN(n1086) );
  XOR2_X2 U896 ( .A(in_b_mac[11]), .B(n1553), .Z(n1072) );
  OAI22_X2 U897 ( .A1(n361), .A2(n1103), .B1(n1068), .B2(n360), .ZN(n1101) );
  XOR2_X2 U898 ( .A(in_b_mac[9]), .B(n1554), .Z(n1068) );
  XNOR2_X2 U900 ( .A(in_b_mac[15]), .B(n230), .ZN(n1089) );
  XOR2_X2 U902 ( .A(n436), .B(in_a_mac[8]), .Z(n1104) );
  OAI22_X2 U904 ( .A1(n361), .A2(n1105), .B1(n1103), .B2(n360), .ZN(n1080) );
  XOR2_X2 U905 ( .A(in_b_mac[10]), .B(n1554), .Z(n1103) );
  XOR2_X2 U909 ( .A(n12), .B(n1109), .Z(n1108) );
  OAI22_X2 U915 ( .A1(n437), .A2(n1113), .B1(n1102), .B2(n814), .ZN(n1074) );
  XOR2_X2 U916 ( .A(in_b_mac[12]), .B(n1553), .Z(n1102) );
  OAI22_X2 U917 ( .A1(n438), .A2(n1111), .B1(n1099), .B2(n721), .ZN(n1076) );
  XOR2_X2 U919 ( .A(in_a_mac[11]), .B(in_a_mac[10]), .Z(n1114) );
  XOR2_X2 U920 ( .A(in_b_mac[14]), .B(n1552), .Z(n1099) );
  XOR2_X2 U921 ( .A(in_b_mac[15]), .B(n1552), .Z(n1111) );
  OAI22_X2 U923 ( .A1(n361), .A2(n1115), .B1(n1105), .B2(n360), .ZN(n1096) );
  XOR2_X2 U924 ( .A(in_b_mac[11]), .B(n1554), .Z(n1105) );
  OAI22_X2 U927 ( .A1(n437), .A2(n1117), .B1(n1113), .B2(n814), .ZN(n1092) );
  XOR2_X2 U928 ( .A(in_b_mac[13]), .B(n1553), .Z(n1113) );
  OAI22_X2 U932 ( .A1(n361), .A2(n368), .B1(n1120), .B2(n360), .ZN(n367) );
  XOR2_X2 U933 ( .A(in_b_mac[14]), .B(n1554), .Z(n368) );
  XOR2_X2 U934 ( .A(U1_C_28_), .B(n12), .Z(n1119) );
  OAI22_X2 U937 ( .A1(n361), .A2(n1120), .B1(n1115), .B2(n360), .ZN(n1107) );
  XOR2_X2 U939 ( .A(in_a_mac[15]), .B(in_a_mac[14]), .Z(n1122) );
  XOR2_X2 U940 ( .A(in_b_mac[12]), .B(n1554), .Z(n1115) );
  XOR2_X2 U941 ( .A(in_b_mac[13]), .B(n1554), .Z(n1120) );
  XNOR2_X2 U942 ( .A(in_a_mac[14]), .B(in_a_mac[13]), .ZN(n361) );
  OAI22_X2 U943 ( .A1(n437), .A2(n1123), .B1(n1117), .B2(n814), .ZN(n1109) );
  XOR2_X2 U944 ( .A(in_b_mac[14]), .B(n1553), .Z(n1117) );
  XOR2_X2 U946 ( .A(in_b_mac[15]), .B(n1553), .Z(n1123) );
  XOR2_X2 U948 ( .A(in_a_mac[13]), .B(in_a_mac[12]), .Z(n1124) );
  OR2_X1 U1158 ( .A1(n443), .A2(n438), .ZN(n720) );
  AND2_X1 U1159 ( .A1(n673), .A2(n672), .ZN(n750) );
  OR2_X1 U1161 ( .A1(n443), .A2(n437), .ZN(n815) );
  AND2_X1 U1162 ( .A1(n798), .A2(n797), .ZN(n861) );
  OR2_X1 U1163 ( .A1(n443), .A2(n361), .ZN(n868) );
  AND2_X1 U1165 ( .A1(n883), .A2(n1502), .ZN(n925) );
  AND2_X1 U1166 ( .A1(n921), .A2(n920), .ZN(n1001) );
  DFF_X2 in_c_mac_reg_30_ ( .D(U6_Z_30), .CK(clk), .Q(U1_C_30_), .QN(n1388) );
  DFF_X2 min_reg_13_ ( .D(U5_Z_13), .CK(clk), .Q(min[13]) );
  DFF_X2 min_reg_12_ ( .D(U5_Z_12), .CK(clk), .Q(min[12]) );
  DFF_X2 min_reg_8_ ( .D(U5_Z_8), .CK(clk), .Q(min[8]) );
  DFF_X2 min_reg_10_ ( .D(U5_Z_10), .CK(clk), .Q(min[10]) );
  DFF_X2 min_reg_9_ ( .D(U5_Z_9), .CK(clk), .Q(min[9]) );
  DFF_X2 min_reg_4_ ( .D(U5_Z_4), .CK(clk), .Q(min[4]) );
  DFF_X2 min_reg_3_ ( .D(U5_Z_3), .CK(clk), .Q(min[3]) );
  DFF_X2 in_c_mac_reg_26_ ( .D(U6_Z_26), .CK(clk), .Q(U1_C_26_) );
  DFF_X2 in_c_mac_reg_31_ ( .D(n424), .CK(clk), .Q(U1_C_31_) );
  DFF_X2 min_reg_11_ ( .D(U5_Z_11), .CK(clk), .Q(min[11]) );
  DFF_X2 min_reg_0_ ( .D(U5_Z_0), .CK(clk), .Q(min[0]) );
  DFF_X2 min_reg_2_ ( .D(U5_Z_2), .CK(clk), .Q(min[2]) );
  DFF_X2 in_c_mac_reg_25_ ( .D(U6_Z_25), .CK(clk), .Q(U1_C_25_), .QN(n18) );
  DFF_X2 in_c_mac_reg_27_ ( .D(U6_Z_27), .CK(clk), .Q(U1_C_27_), .QN(n12) );
  DFF_X2 in_c_mac_reg_0_ ( .D(U6_Z_0), .CK(clk), .Q(U1_C_0_), .QN(n490) );
  DFF_X2 in_c_mac_reg_1_ ( .D(U6_Z_1), .CK(clk), .Q(U1_C_1_) );
  DFF_X2 in_c_mac_reg_2_ ( .D(U6_Z_2), .CK(clk), .Q(U1_C_2_), .QN(n512) );
  DFF_X2 in_c_mac_reg_3_ ( .D(U6_Z_3), .CK(clk), .Q(U1_C_3_) );
  DFF_X2 in_c_mac_reg_4_ ( .D(U6_Z_4), .CK(clk), .Q(U1_C_4_) );
  DFF_X2 in_c_mac_reg_5_ ( .D(U6_Z_5), .CK(clk), .Q(U1_C_5_) );
  DFF_X2 in_c_mac_reg_6_ ( .D(U6_Z_6), .CK(clk), .Q(U1_C_6_) );
  DFF_X2 in_c_mac_reg_7_ ( .D(U6_Z_7), .CK(clk), .Q(U1_C_7_) );
  DFF_X2 in_c_mac_reg_8_ ( .D(U6_Z_8), .CK(clk), .Q(U1_C_8_) );
  DFF_X2 in_c_mac_reg_9_ ( .D(U6_Z_9), .CK(clk), .Q(U1_C_9_) );
  DFF_X2 in_c_mac_reg_12_ ( .D(U6_Z_12), .CK(clk), .Q(U1_C_12_), .QN(n467) );
  DFF_X2 in_c_mac_reg_10_ ( .D(U6_Z_10), .CK(clk), .Q(U1_C_10_), .QN(n476) );
  DFF_X2 in_c_mac_reg_11_ ( .D(U6_Z_11), .CK(clk), .Q(U1_C_11_) );
  DFF_X2 in_c_mac_reg_13_ ( .D(U6_Z_13), .CK(clk), .Q(U1_C_13_) );
  DFF_X2 in_c_mac_reg_14_ ( .D(U6_Z_14), .CK(clk), .Q(U1_C_14_), .QN(n617) );
  DFF_X2 in_c_mac_reg_15_ ( .D(U6_Z_15), .CK(clk), .Q(U1_C_15_) );
  DFF_X2 in_c_mac_reg_16_ ( .D(U6_Z_16), .CK(clk), .Q(U1_C_16_) );
  DFF_X2 in_c_mac_reg_18_ ( .D(U6_Z_18), .CK(clk), .Q(U1_C_18_) );
  DFF_X2 in_c_mac_reg_20_ ( .D(U6_Z_20), .CK(clk), .Q(U1_C_20_) );
  DFF_X2 in_c_mac_reg_22_ ( .D(U6_Z_22), .CK(clk), .Q(U1_C_22_) );
  DFF_X2 in_c_mac_reg_24_ ( .D(U6_Z_24), .CK(clk), .Q(U1_C_24_) );
  DFF_X2 in_c_mac_reg_28_ ( .D(U6_Z_28), .CK(clk), .Q(U1_C_28_) );
  DFF_X2 in_c_mac_reg_17_ ( .D(U6_Z_17), .CK(clk), .Q(U1_C_17_), .QN(n65) );
  DFF_X2 in_c_mac_reg_19_ ( .D(U6_Z_19), .CK(clk), .Q(n593), .QN(n52) );
  DFF_X2 in_c_mac_reg_21_ ( .D(U6_Z_21), .CK(clk), .Q(U1_C_21_), .QN(n41) );
  DFF_X2 in_c_mac_reg_23_ ( .D(U6_Z_23), .CK(clk), .Q(U1_C_23_), .QN(n29) );
  DFF_X2 in_c_mac_reg_29_ ( .D(U6_Z_29), .CK(clk), .Q(n1367), .QN(n4) );
  DFF_X2 min_reg_14_ ( .D(U5_Z_14), .CK(clk), .Q(min[14]) );
  DFF_X2 min_reg_7_ ( .D(U5_Z_7), .CK(clk), .Q(min[7]) );
  DFF_X2 min_reg_6_ ( .D(U5_Z_6), .CK(clk), .Q(min[6]) );
  DFF_X2 min_reg_5_ ( .D(U5_Z_5), .CK(clk), .Q(min[5]) );
  DFF_X2 min_reg_1_ ( .D(U5_Z_1), .CK(clk), .Q(min[1]) );
  INV_X4 U8 ( .A(n433), .ZN(n434) );
  OAI21_X2 U10 ( .B1(n850), .B2(n1491), .A(n839), .ZN(n902) );
  NAND2_X2 U11 ( .A1(n1383), .A2(n180), .ZN(n181) );
  NAND2_X2 U13 ( .A1(n179), .A2(n1387), .ZN(n182) );
  NAND2_X2 U14 ( .A1(n181), .A2(n182), .ZN(n1381) );
  INV_X1 U15 ( .A(n1383), .ZN(n179) );
  INV_X4 U16 ( .A(n1387), .ZN(n180) );
  INV_X1 U17 ( .A(n241), .ZN(n857) );
  NOR2_X1 U18 ( .A1(n241), .A2(n851), .ZN(n855) );
  NOR2_X4 U19 ( .A1(n1425), .A2(n1314), .ZN(n1315) );
  NAND2_X2 U20 ( .A1(n431), .A2(n445), .ZN(n1445) );
  NOR2_X2 U21 ( .A1(n1409), .A2(n1255), .ZN(n1264) );
  NAND2_X2 U22 ( .A1(n563), .A2(U1_C_5_), .ZN(n781) );
  NOR2_X2 U23 ( .A1(n1482), .A2(n1480), .ZN(n1157) );
  OAI21_X2 U24 ( .B1(n1090), .B2(n1472), .A(n1073), .ZN(n1477) );
  NAND2_X2 U25 ( .A1(n555), .A2(n556), .ZN(n577) );
  INV_X4 U26 ( .A(in_a_mac[1]), .ZN(n433) );
  NAND2_X2 U27 ( .A1(n569), .A2(n214), .ZN(n185) );
  NAND2_X2 U28 ( .A1(n183), .A2(n184), .ZN(n186) );
  NAND2_X2 U33 ( .A1(n185), .A2(n186), .ZN(n393) );
  INV_X4 U34 ( .A(n569), .ZN(n183) );
  INV_X4 U38 ( .A(n214), .ZN(n184) );
  NAND2_X2 U39 ( .A1(n951), .A2(n950), .ZN(n189) );
  NAND2_X2 U40 ( .A1(n187), .A2(n188), .ZN(n190) );
  NAND2_X2 U46 ( .A1(n189), .A2(n190), .ZN(n369) );
  INV_X4 U47 ( .A(n951), .ZN(n187) );
  INV_X4 U49 ( .A(n950), .ZN(n188) );
  NAND2_X2 U50 ( .A1(n414), .A2(n511), .ZN(n192) );
  NAND2_X2 U52 ( .A1(n191), .A2(n515), .ZN(n193) );
  NAND2_X2 U53 ( .A1(n192), .A2(n193), .ZN(n510) );
  INV_X4 U55 ( .A(n414), .ZN(n191) );
  NAND2_X1 U56 ( .A1(n443), .A2(n235), .ZN(n511) );
  NAND2_X2 U58 ( .A1(n338), .A2(n562), .ZN(n195) );
  NAND2_X2 U59 ( .A1(n194), .A2(n558), .ZN(n196) );
  NAND2_X2 U61 ( .A1(n195), .A2(n196), .ZN(n569) );
  INV_X4 U62 ( .A(n338), .ZN(n194) );
  NAND2_X2 U63 ( .A1(n566), .A2(n782), .ZN(n198) );
  NAND2_X2 U64 ( .A1(n197), .A2(n786), .ZN(n199) );
  NAND2_X2 U65 ( .A1(n198), .A2(n199), .ZN(n767) );
  INV_X4 U66 ( .A(n566), .ZN(n197) );
  NAND2_X2 U67 ( .A1(in_a_mac[2]), .A2(n433), .ZN(n201) );
  NAND2_X2 U68 ( .A1(n200), .A2(in_a_mac[1]), .ZN(n202) );
  NAND2_X2 U69 ( .A1(n201), .A2(n202), .ZN(n416) );
  INV_X4 U70 ( .A(in_a_mac[2]), .ZN(n200) );
  NAND2_X2 U71 ( .A1(n1392), .A2(n322), .ZN(n205) );
  NAND2_X2 U72 ( .A1(n203), .A2(n204), .ZN(n206) );
  NAND2_X2 U73 ( .A1(n205), .A2(n206), .ZN(n321) );
  INV_X4 U74 ( .A(n1392), .ZN(n203) );
  INV_X4 U75 ( .A(n322), .ZN(n204) );
  NAND2_X2 U76 ( .A1(n413), .A2(n375), .ZN(n211) );
  NAND2_X2 U77 ( .A1(n207), .A2(n210), .ZN(n213) );
  NAND2_X2 U78 ( .A1(n211), .A2(n213), .ZN(n538) );
  INV_X4 U79 ( .A(n413), .ZN(n207) );
  INV_X4 U80 ( .A(n375), .ZN(n210) );
  AND2_X4 U81 ( .A1(n443), .A2(n542), .ZN(n375) );
  OAI21_X2 U82 ( .B1(n577), .B2(n576), .A(n575), .ZN(n578) );
  INV_X2 U83 ( .A(n1380), .ZN(n1375) );
  NOR2_X2 U84 ( .A1(n754), .A2(n751), .ZN(n1458) );
  AOI21_X2 U85 ( .B1(n815), .B2(n814), .A(n1553), .ZN(n709) );
  INV_X4 U86 ( .A(in_b_mac[5]), .ZN(n251) );
  INV_X4 U87 ( .A(n1476), .ZN(n301) );
  NAND2_X2 U88 ( .A1(n438), .A2(n1114), .ZN(n721) );
  OAI21_X2 U89 ( .B1(n1547), .B2(n1549), .A(n810), .ZN(n740) );
  INV_X4 U90 ( .A(in_b_mac[4]), .ZN(n332) );
  INV_X4 U91 ( .A(n428), .ZN(n352) );
  OAI21_X2 U92 ( .B1(n732), .B2(n731), .A(n729), .ZN(n799) );
  AOI21_X2 U93 ( .B1(n698), .B2(n700), .A(n701), .ZN(n776) );
  AOI21_X2 U94 ( .B1(n789), .B2(n1242), .A(n907), .ZN(n842) );
  NAND2_X2 U95 ( .A1(n437), .A2(n1124), .ZN(n814) );
  NAND2_X2 U96 ( .A1(n361), .A2(n1122), .ZN(n360) );
  AOI21_X2 U97 ( .B1(n624), .B2(n623), .A(n621), .ZN(n688) );
  NAND2_X2 U98 ( .A1(n578), .A2(n579), .ZN(n753) );
  OAI22_X2 U99 ( .A1(n1358), .A2(n1357), .B1(n1356), .B2(n1355), .ZN(n1438) );
  NOR2_X2 U100 ( .A1(n1375), .A2(n1376), .ZN(n1377) );
  INV_X1 U101 ( .A(n314), .ZN(n312) );
  INV_X2 U102 ( .A(n780), .ZN(n850) );
  INV_X4 U103 ( .A(n1493), .ZN(n834) );
  XNOR2_X1 U104 ( .A(n668), .B(n315), .ZN(n564) );
  INV_X2 U105 ( .A(n1428), .ZN(n1330) );
  INV_X2 U106 ( .A(n1344), .ZN(n326) );
  INV_X2 U107 ( .A(n1191), .ZN(n298) );
  XNOR2_X1 U108 ( .A(n563), .B(U1_C_5_), .ZN(n214) );
  INV_X4 U109 ( .A(n1233), .ZN(n314) );
  INV_X4 U110 ( .A(in_b_mac[0]), .ZN(n444) );
  INV_X4 U111 ( .A(n444), .ZN(n443) );
  OAI22_X1 U112 ( .A1(n1504), .A2(n1503), .B1(n1156), .B2(n1155), .ZN(n1160)
         );
  INV_X4 U113 ( .A(in_a_mac[5]), .ZN(n668) );
  OAI22_X1 U114 ( .A1(n857), .A2(n856), .B1(n855), .B2(n853), .ZN(n904) );
  XNOR2_X2 U115 ( .A(n1366), .B(n300), .ZN(n215) );
  XOR2_X2 U116 ( .A(n823), .B(n404), .Z(n216) );
  AND2_X4 U117 ( .A1(n569), .A2(n568), .ZN(n218) );
  OAI21_X1 U118 ( .B1(n218), .B2(n214), .A(n571), .ZN(n752) );
  INV_X4 U119 ( .A(n417), .ZN(n438) );
  XOR2_X1 U120 ( .A(in_a_mac[10]), .B(n436), .Z(n417) );
  INV_X4 U121 ( .A(n421), .ZN(n437) );
  XNOR2_X2 U122 ( .A(n1441), .B(n923), .ZN(n219) );
  NOR2_X2 U123 ( .A1(n822), .A2(n1215), .ZN(n220) );
  XNOR2_X2 U124 ( .A(n1426), .B(n334), .ZN(n221) );
  XNOR2_X2 U125 ( .A(n1273), .B(n959), .ZN(n222) );
  OAI22_X1 U126 ( .A1(n438), .A2(n984), .B1(n948), .B2(n721), .ZN(n982) );
  XNOR2_X2 U127 ( .A(n1287), .B(n992), .ZN(n223) );
  AND2_X4 U128 ( .A1(n1121), .A2(n633), .ZN(n224) );
  NOR2_X4 U129 ( .A1(n1428), .A2(n1429), .ZN(n1328) );
  INV_X1 U130 ( .A(n1482), .ZN(n225) );
  INV_X4 U131 ( .A(n1159), .ZN(n1482) );
  NOR2_X2 U133 ( .A1(n1436), .A2(n1434), .ZN(n1350) );
  INV_X1 U134 ( .A(n1436), .ZN(n292) );
  INV_X1 U135 ( .A(n1165), .ZN(n337) );
  INV_X1 U136 ( .A(n1425), .ZN(n333) );
  NOR2_X2 U137 ( .A1(n314), .A2(n1228), .ZN(n1232) );
  NOR2_X2 U138 ( .A1(n1395), .A2(n1393), .ZN(n1204) );
  NOR2_X4 U139 ( .A1(n1165), .A2(n1483), .ZN(n1175) );
  NAND3_X1 U140 ( .A1(n759), .A2(n579), .A3(n578), .ZN(n763) );
  OAI22_X2 U141 ( .A1(n1487), .A2(n1190), .B1(n1489), .B2(n1191), .ZN(n226) );
  INV_X4 U142 ( .A(n226), .ZN(n1395) );
  OAI22_X2 U143 ( .A1(n1363), .A2(n1364), .B1(n1365), .B2(n1438), .ZN(n1380)
         );
  OAI22_X2 U144 ( .A1(n1315), .A2(n1423), .B1(n1424), .B2(n1316), .ZN(n1428)
         );
  OAI22_X2 U145 ( .A1(n1431), .A2(n1343), .B1(n1432), .B2(n1344), .ZN(n1351)
         );
  OAI22_X2 U146 ( .A1(n1377), .A2(n1378), .B1(n1380), .B2(n1379), .ZN(n1386)
         );
  OAI22_X2 U147 ( .A1(n1157), .A2(n1479), .B1(n1159), .B2(n1158), .ZN(n1485)
         );
  OAI22_X2 U148 ( .A1(n1175), .A2(n1484), .B1(n1176), .B2(n1485), .ZN(n1191)
         );
  OAI22_X2 U149 ( .A1(n961), .A2(n1467), .B1(n969), .B2(n968), .ZN(n1471) );
  XNOR2_X2 U150 ( .A(n433), .B(n315), .ZN(n496) );
  INV_X4 U151 ( .A(in_b_mac[1]), .ZN(n315) );
  XNOR2_X2 U152 ( .A(n567), .B(n768), .ZN(n755) );
  OAI22_X1 U153 ( .A1(n562), .A2(n561), .B1(n560), .B2(n329), .ZN(n773) );
  INV_X4 U154 ( .A(n439), .ZN(n440) );
  INV_X1 U155 ( .A(n613), .ZN(n439) );
  XNOR2_X2 U156 ( .A(n678), .B(n661), .ZN(n372) );
  INV_X2 U157 ( .A(n661), .ZN(n1548) );
  OAI21_X2 U158 ( .B1(n664), .B2(n1550), .A(n230), .ZN(n661) );
  INV_X4 U159 ( .A(n550), .ZN(n548) );
  NAND2_X2 U160 ( .A1(n761), .A2(n763), .ZN(n227) );
  NAND2_X2 U161 ( .A1(n761), .A2(n763), .ZN(n1493) );
  NAND2_X2 U162 ( .A1(n275), .A2(n1475), .ZN(n309) );
  INV_X2 U163 ( .A(n1477), .ZN(n275) );
  OAI22_X1 U164 ( .A1(n1127), .A2(n1126), .B1(n1125), .B2(n1118), .ZN(n1140)
         );
  INV_X1 U165 ( .A(n292), .ZN(n228) );
  NAND2_X1 U166 ( .A1(n570), .A2(n183), .ZN(n571) );
  XNOR2_X2 U167 ( .A(n807), .B(n792), .ZN(n853) );
  XOR2_X1 U168 ( .A(n790), .B(n788), .Z(n807) );
  OAI22_X1 U169 ( .A1(n491), .A2(n490), .B1(n489), .B2(n433), .ZN(n492) );
  INV_X1 U170 ( .A(n436), .ZN(n229) );
  INV_X4 U171 ( .A(n229), .ZN(n230) );
  INV_X4 U172 ( .A(n435), .ZN(n436) );
  XOR2_X1 U173 ( .A(n428), .B(n319), .Z(n565) );
  INV_X1 U174 ( .A(n758), .ZN(n231) );
  INV_X4 U175 ( .A(n231), .ZN(n232) );
  INV_X1 U176 ( .A(n529), .ZN(n233) );
  INV_X4 U177 ( .A(n233), .ZN(n234) );
  XNOR2_X2 U178 ( .A(n241), .B(n853), .ZN(n831) );
  XNOR2_X2 U179 ( .A(n433), .B(n319), .ZN(n525) );
  NAND2_X4 U180 ( .A1(in_a_mac[1]), .A2(n717), .ZN(n716) );
  INV_X16 U181 ( .A(in_a_mac[0]), .ZN(n717) );
  NOR2_X1 U182 ( .A1(n493), .A2(n492), .ZN(n495) );
  INV_X1 U183 ( .A(n498), .ZN(n494) );
  XNOR2_X2 U184 ( .A(in_a_mac[2]), .B(n427), .ZN(n461) );
  INV_X1 U185 ( .A(n432), .ZN(n235) );
  INV_X4 U186 ( .A(n235), .ZN(n236) );
  INV_X4 U187 ( .A(n416), .ZN(n432) );
  NOR2_X2 U188 ( .A1(n541), .A2(n1445), .ZN(n331) );
  XNOR2_X2 U189 ( .A(in_a_mac[5]), .B(n443), .ZN(n541) );
  XNOR2_X2 U190 ( .A(n237), .B(n934), .ZN(n1495) );
  XNOR2_X2 U191 ( .A(n936), .B(n917), .ZN(n237) );
  INV_X2 U192 ( .A(n934), .ZN(n915) );
  OAI22_X1 U193 ( .A1(n901), .A2(n894), .B1(n891), .B2(n307), .ZN(n934) );
  OAI22_X1 U194 ( .A1(n716), .A2(n443), .B1(n717), .B2(n496), .ZN(n252) );
  XOR2_X1 U195 ( .A(n427), .B(in_b_mac[6]), .Z(n238) );
  XOR2_X1 U196 ( .A(n427), .B(in_b_mac[6]), .Z(n659) );
  INV_X4 U197 ( .A(in_a_mac[3]), .ZN(n427) );
  INV_X1 U198 ( .A(n573), .ZN(n239) );
  INV_X4 U199 ( .A(n239), .ZN(n240) );
  XNOR2_X2 U200 ( .A(n391), .B(n894), .ZN(n241) );
  INV_X4 U201 ( .A(in_b_mac[3]), .ZN(n319) );
  XNOR2_X1 U202 ( .A(in_a_mac[8]), .B(in_a_mac[7]), .ZN(n613) );
  INV_X4 U203 ( .A(in_a_mac[7]), .ZN(n1551) );
  OAI22_X1 U204 ( .A1(n546), .A2(n717), .B1(n525), .B2(n716), .ZN(n246) );
  INV_X2 U205 ( .A(n1395), .ZN(n335) );
  XNOR2_X2 U206 ( .A(n251), .B(n433), .ZN(n559) );
  NAND2_X2 U207 ( .A1(n544), .A2(in_a_mac[5]), .ZN(n561) );
  NAND2_X2 U208 ( .A1(n432), .A2(n461), .ZN(n253) );
  OAI22_X1 U209 ( .A1(n945), .A2(n1442), .B1(n944), .B2(n430), .ZN(n911) );
  OAI22_X1 U210 ( .A1(n860), .A2(n1442), .B1(n945), .B2(n430), .ZN(n898) );
  OAI22_X1 U211 ( .A1(n1041), .A2(n1442), .B1(n1056), .B2(n430), .ZN(n1037) );
  OAI22_X1 U212 ( .A1(n976), .A2(n430), .B1(n944), .B2(n1442), .ZN(n610) );
  OAI22_X1 U213 ( .A1(n1016), .A2(n430), .B1(n976), .B2(n1442), .ZN(n599) );
  OAI22_X1 U214 ( .A1(n1041), .A2(n430), .B1(n1016), .B2(n1442), .ZN(n1259) );
  OAI22_X1 U215 ( .A1(n726), .A2(n430), .B1(n692), .B2(n1442), .ZN(n981) );
  OAI22_X1 U216 ( .A1(n760), .A2(n430), .B1(n726), .B2(n1442), .ZN(n1128) );
  OAI22_X1 U217 ( .A1(n820), .A2(n430), .B1(n760), .B2(n1442), .ZN(n751) );
  OAI22_X1 U218 ( .A1(n830), .A2(n430), .B1(n820), .B2(n1442), .ZN(n455) );
  OAI22_X1 U219 ( .A1(n860), .A2(n430), .B1(n830), .B2(n1442), .ZN(n446) );
  AND2_X1 U220 ( .A1(n719), .A2(n1442), .ZN(n395) );
  NAND2_X2 U221 ( .A1(n432), .A2(n461), .ZN(n254) );
  XNOR2_X2 U222 ( .A(n867), .B(n866), .ZN(n380) );
  INV_X4 U223 ( .A(n753), .ZN(n758) );
  INV_X1 U224 ( .A(n950), .ZN(n260) );
  INV_X1 U225 ( .A(n532), .ZN(n261) );
  INV_X4 U226 ( .A(n261), .ZN(n262) );
  NOR2_X1 U227 ( .A1(n955), .A2(n953), .ZN(n263) );
  NOR2_X1 U228 ( .A1(n325), .A2(n1405), .ZN(n265) );
  INV_X1 U229 ( .A(n553), .ZN(n266) );
  XNOR2_X2 U230 ( .A(n778), .B(n772), .ZN(n567) );
  INV_X1 U231 ( .A(n253), .ZN(n267) );
  INV_X4 U232 ( .A(n267), .ZN(n268) );
  INV_X1 U233 ( .A(n712), .ZN(n270) );
  OAI22_X2 U234 ( .A1(n546), .A2(n717), .B1(n525), .B2(n716), .ZN(n287) );
  INV_X2 U235 ( .A(n1491), .ZN(n1492) );
  INV_X1 U236 ( .A(n520), .ZN(n271) );
  INV_X1 U237 ( .A(n523), .ZN(n520) );
  INV_X1 U238 ( .A(n1445), .ZN(n272) );
  INV_X2 U239 ( .A(n272), .ZN(n273) );
  NOR2_X2 U240 ( .A1(n282), .A2(n208), .ZN(n424) );
  INV_X4 U241 ( .A(n275), .ZN(n276) );
  OAI22_X2 U242 ( .A1(U1_C_4_), .A2(n246), .B1(n375), .B2(n547), .ZN(n568) );
  INV_X1 U243 ( .A(n916), .ZN(n277) );
  INV_X1 U244 ( .A(n936), .ZN(n916) );
  INV_X1 U245 ( .A(n548), .ZN(n278) );
  NAND2_X1 U246 ( .A1(n613), .A2(n1104), .ZN(n280) );
  NAND2_X2 U247 ( .A1(n613), .A2(n1104), .ZN(n642) );
  INV_X1 U248 ( .A(n1498), .ZN(n1499) );
  XNOR2_X2 U249 ( .A(n828), .B(U1_C_6_), .ZN(n411) );
  AOI21_X2 U250 ( .B1(n656), .B2(n657), .A(n1543), .ZN(n281) );
  AOI21_X2 U251 ( .B1(n720), .B2(n721), .A(n1552), .ZN(n657) );
  AOI21_X2 U252 ( .B1(n656), .B2(n657), .A(n1543), .ZN(n647) );
  INV_X2 U253 ( .A(n415), .ZN(n282) );
  XNOR2_X2 U254 ( .A(n538), .B(n540), .ZN(n527) );
  INV_X2 U255 ( .A(n535), .ZN(n540) );
  INV_X2 U256 ( .A(n284), .ZN(n1291) );
  OAI22_X1 U257 ( .A1(n1411), .A2(n1279), .B1(n1278), .B2(n1277), .ZN(n284) );
  AOI21_X4 U258 ( .B1(n1500), .B2(n1501), .A(n1498), .ZN(n955) );
  OAI21_X4 U259 ( .B1(n914), .B2(n1495), .A(n906), .ZN(n1500) );
  NOR2_X4 U260 ( .A1(n1496), .A2(n1497), .ZN(n914) );
  INV_X1 U261 ( .A(n1500), .ZN(n285) );
  INV_X4 U262 ( .A(n285), .ZN(n286) );
  INV_X1 U263 ( .A(n1303), .ZN(n288) );
  INV_X1 U264 ( .A(n1291), .ZN(n289) );
  INV_X1 U265 ( .A(n1330), .ZN(n290) );
  INV_X1 U266 ( .A(n1220), .ZN(n291) );
  INV_X2 U267 ( .A(n1271), .ZN(n1411) );
  OAI22_X1 U268 ( .A1(n313), .A2(n1247), .B1(n265), .B2(n1245), .ZN(n293) );
  INV_X1 U269 ( .A(n1365), .ZN(n294) );
  NOR2_X2 U270 ( .A1(n326), .A2(n1338), .ZN(n1343) );
  INV_X1 U271 ( .A(n834), .ZN(n295) );
  NOR2_X1 U272 ( .A1(n396), .A2(n415), .ZN(U5_Z_14) );
  INV_X4 U273 ( .A(n552), .ZN(n553) );
  INV_X1 U274 ( .A(n1191), .ZN(n1490) );
  NOR2_X2 U275 ( .A1(n298), .A2(n1189), .ZN(n1190) );
  INV_X4 U276 ( .A(n1490), .ZN(n429) );
  INV_X1 U277 ( .A(n577), .ZN(n296) );
  INV_X4 U278 ( .A(n296), .ZN(n297) );
  NOR2_X2 U279 ( .A1(n1416), .A2(n1285), .ZN(n1290) );
  INV_X1 U280 ( .A(n225), .ZN(n299) );
  INV_X1 U281 ( .A(n1380), .ZN(n300) );
  NOR2_X2 U282 ( .A1(n325), .A2(n1405), .ZN(n1246) );
  INV_X4 U283 ( .A(n1351), .ZN(n1436) );
  INV_X4 U284 ( .A(n333), .ZN(n334) );
  NAND2_X2 U285 ( .A1(n302), .A2(n301), .ZN(n310) );
  NAND2_X2 U286 ( .A1(n1477), .A2(n1140), .ZN(n302) );
  XNOR2_X2 U287 ( .A(n781), .B(n426), .ZN(n566) );
  XOR2_X1 U288 ( .A(n352), .B(in_b_mac[4]), .Z(n819) );
  XOR2_X1 U289 ( .A(n352), .B(in_b_mac[5]), .Z(n824) );
  OAI22_X1 U290 ( .A1(n778), .A2(n773), .B1(n771), .B2(n772), .ZN(n1494) );
  NAND2_X1 U291 ( .A1(n329), .A2(n561), .ZN(n305) );
  NAND2_X2 U292 ( .A1(n303), .A2(n304), .ZN(n306) );
  NAND2_X2 U293 ( .A1(n305), .A2(n306), .ZN(n338) );
  INV_X1 U294 ( .A(n329), .ZN(n303) );
  INV_X1 U295 ( .A(n561), .ZN(n304) );
  NOR2_X2 U296 ( .A1(n330), .A2(n331), .ZN(n329) );
  XNOR2_X2 U297 ( .A(n818), .B(U1_C_7_), .ZN(n307) );
  INV_X4 U298 ( .A(n307), .ZN(n882) );
  INV_X4 U299 ( .A(n321), .ZN(n415) );
  INV_X1 U300 ( .A(n1383), .ZN(n308) );
  NAND2_X2 U301 ( .A1(n309), .A2(n310), .ZN(n1159) );
  INV_X1 U302 ( .A(n1344), .ZN(n311) );
  INV_X2 U303 ( .A(n325), .ZN(n313) );
  INV_X1 U304 ( .A(n1439), .ZN(n1363) );
  NOR2_X2 U305 ( .A1(n431), .A2(n564), .ZN(n330) );
  OAI22_X2 U306 ( .A1(n559), .A2(n717), .B1(n546), .B2(n716), .ZN(n563) );
  OAI22_X2 U307 ( .A1(n443), .A2(n716), .B1(n717), .B2(n496), .ZN(n487) );
  INV_X1 U308 ( .A(n312), .ZN(n1403) );
  INV_X1 U309 ( .A(in_b_mac[2]), .ZN(n316) );
  INV_X4 U310 ( .A(n316), .ZN(n317) );
  NAND2_X1 U311 ( .A1(n443), .A2(n454), .ZN(n615) );
  XOR2_X1 U312 ( .A(n1554), .B(n443), .Z(n872) );
  NAND2_X1 U313 ( .A1(n443), .A2(n421), .ZN(n468) );
  XOR2_X1 U314 ( .A(n1553), .B(n443), .Z(n813) );
  AND2_X1 U315 ( .A1(n443), .A2(n439), .ZN(n402) );
  NAND2_X1 U316 ( .A1(n443), .A2(n417), .ZN(n680) );
  NOR2_X1 U317 ( .A1(n443), .A2(n613), .ZN(n664) );
  NAND2_X1 U318 ( .A1(in_a_mac[0]), .A2(n443), .ZN(n491) );
  XOR2_X1 U319 ( .A(n1551), .B(n443), .Z(n596) );
  XNOR2_X1 U320 ( .A(n443), .B(n428), .ZN(n505) );
  XNOR2_X1 U321 ( .A(in_b_mac[3]), .B(n436), .ZN(n722) );
  XOR2_X1 U322 ( .A(in_b_mac[3]), .B(n1551), .Z(n665) );
  INV_X8 U323 ( .A(n419), .ZN(n430) );
  INV_X2 U324 ( .A(n737), .ZN(n738) );
  INV_X1 U325 ( .A(n1397), .ZN(n1220) );
  OAI22_X1 U326 ( .A1(U1_C_2_), .A2(n516), .B1(n515), .B2(n514), .ZN(n530) );
  INV_X1 U327 ( .A(n431), .ZN(n542) );
  INV_X4 U328 ( .A(n1485), .ZN(n1165) );
  XOR2_X2 U330 ( .A(in_a_mac[4]), .B(in_a_mac[5]), .Z(n445) );
  AND2_X4 U331 ( .A1(n434), .A2(n717), .ZN(n318) );
  NAND2_X1 U332 ( .A1(U1_C_7_), .A2(n818), .ZN(n736) );
  INV_X4 U333 ( .A(n319), .ZN(n320) );
  XNOR2_X1 U334 ( .A(in_b_mac[12]), .B(n434), .ZN(n746) );
  XNOR2_X1 U335 ( .A(in_b_mac[10]), .B(n434), .ZN(n696) );
  XNOR2_X1 U336 ( .A(in_b_mac[11]), .B(n434), .ZN(n747) );
  XNOR2_X1 U337 ( .A(in_b_mac[9]), .B(n434), .ZN(n660) );
  XOR2_X2 U338 ( .A(U1_C_31_), .B(n1391), .Z(n322) );
  INV_X1 U339 ( .A(n1496), .ZN(n323) );
  INV_X4 U340 ( .A(n323), .ZN(n324) );
  INV_X4 U341 ( .A(n1316), .ZN(n1425) );
  INV_X4 U342 ( .A(n1248), .ZN(n325) );
  NOR2_X2 U343 ( .A1(n955), .A2(n953), .ZN(n1467) );
  INV_X1 U344 ( .A(n1409), .ZN(n327) );
  INV_X4 U345 ( .A(n327), .ZN(n328) );
  XNOR2_X2 U346 ( .A(n433), .B(n332), .ZN(n546) );
  XNOR2_X1 U347 ( .A(in_b_mac[13]), .B(n434), .ZN(n817) );
  XNOR2_X1 U348 ( .A(in_b_mac[15]), .B(n434), .ZN(n896) );
  XNOR2_X1 U349 ( .A(in_b_mac[14]), .B(n434), .ZN(n833) );
  OAI22_X1 U351 ( .A1(n833), .A2(n717), .B1(n817), .B2(n716), .ZN(n622) );
  OAI22_X1 U352 ( .A1(n896), .A2(n717), .B1(n833), .B2(n716), .ZN(n1444) );
  XOR2_X1 U353 ( .A(n668), .B(in_b_mac[15]), .Z(n588) );
  XOR2_X1 U355 ( .A(n668), .B(in_b_mac[11]), .Z(n1446) );
  XOR2_X1 U356 ( .A(n668), .B(in_b_mac[12]), .Z(n1447) );
  XOR2_X1 U357 ( .A(n668), .B(in_b_mac[10]), .Z(n450) );
  XOR2_X1 U358 ( .A(n668), .B(in_b_mac[8]), .Z(n471) );
  XOR2_X1 U359 ( .A(n668), .B(in_b_mac[9]), .Z(n470) );
  XOR2_X1 U360 ( .A(n668), .B(in_b_mac[7]), .Z(n472) );
  XOR2_X1 U361 ( .A(n668), .B(in_b_mac[6]), .Z(n669) );
  XOR2_X1 U362 ( .A(n668), .B(in_b_mac[5]), .Z(n687) );
  XOR2_X1 U363 ( .A(n668), .B(in_b_mac[4]), .Z(n685) );
  XOR2_X1 U364 ( .A(n668), .B(in_b_mac[3]), .Z(n727) );
  XOR2_X1 U365 ( .A(n668), .B(in_b_mac[2]), .Z(n723) );
  OAI22_X1 U366 ( .A1(n236), .A2(n545), .B1(n526), .B2(n253), .ZN(n539) );
  INV_X4 U367 ( .A(n335), .ZN(n336) );
  XOR2_X1 U368 ( .A(n580), .B(n232), .Z(n581) );
  NAND2_X2 U369 ( .A1(n577), .A2(n576), .ZN(n579) );
  OAI21_X4 U370 ( .B1(n758), .B2(n759), .A(n755), .ZN(n761) );
  OAI21_X2 U371 ( .B1(U1_C_3_), .B2(n507), .A(n535), .ZN(n518) );
  OAI22_X2 U372 ( .A1(n525), .A2(n717), .B1(n506), .B2(n716), .ZN(n507) );
  INV_X8 U373 ( .A(n418), .ZN(n431) );
  OAI21_X2 U374 ( .B1(n709), .B2(n811), .A(n710), .ZN(n810) );
  NOR2_X2 U375 ( .A1(n805), .A2(n806), .ZN(n1451) );
  INV_X4 U376 ( .A(in_a_mac[11]), .ZN(n1552) );
  XOR2_X1 U377 ( .A(n380), .B(n875), .Z(n917) );
  AND2_X4 U378 ( .A1(n443), .A2(n718), .ZN(n385) );
  OAI21_X2 U379 ( .B1(n505), .B2(n253), .A(n504), .ZN(n523) );
  XNOR2_X2 U380 ( .A(n346), .B(n748), .ZN(n938) );
  XNOR2_X2 U381 ( .A(n1537), .B(n344), .ZN(n343) );
  INV_X4 U382 ( .A(n558), .ZN(n562) );
  AND2_X4 U383 ( .A1(n561), .A2(n562), .ZN(n560) );
  INV_X1 U384 ( .A(n1126), .ZN(n339) );
  INV_X1 U385 ( .A(n1106), .ZN(n1127) );
  INV_X1 U386 ( .A(n890), .ZN(n1509) );
  AOI21_X1 U387 ( .B1(n841), .B2(n842), .A(n840), .ZN(n884) );
  NOR2_X1 U388 ( .A1(n842), .A2(n841), .ZN(n1243) );
  NAND2_X1 U389 ( .A1(n542), .A2(n444), .ZN(n543) );
  XNOR2_X2 U390 ( .A(n345), .B(n646), .ZN(n1141) );
  XOR2_X2 U391 ( .A(n1132), .B(n647), .Z(n345) );
  INV_X1 U392 ( .A(n1043), .ZN(n342) );
  INV_X1 U394 ( .A(n1017), .ZN(n1044) );
  NOR2_X1 U395 ( .A1(n1017), .A2(n342), .ZN(n1019) );
  INV_X1 U396 ( .A(n899), .ZN(n1513) );
  XOR2_X1 U397 ( .A(n442), .B(in_a_mac[5]), .Z(n627) );
  XOR2_X1 U398 ( .A(n441), .B(in_a_mac[5]), .Z(n602) );
  XOR2_X2 U399 ( .A(in_a_mac[6]), .B(in_a_mac[5]), .Z(n419) );
  AND2_X4 U400 ( .A1(n1163), .A2(n1164), .ZN(n1161) );
  NOR2_X2 U402 ( .A1(n339), .A2(n1106), .ZN(n1118) );
  XOR2_X1 U403 ( .A(n294), .B(n388), .Z(n242) );
  XNOR2_X1 U404 ( .A(n707), .B(n676), .ZN(n675) );
  NOR2_X1 U405 ( .A1(n656), .A2(n657), .ZN(n1464) );
  XNOR2_X2 U406 ( .A(n729), .B(n341), .ZN(n340) );
  XNOR2_X1 U407 ( .A(n731), .B(n732), .ZN(n341) );
  INV_X1 U408 ( .A(n777), .ZN(n383) );
  AOI21_X1 U409 ( .B1(n769), .B2(n220), .A(n766), .ZN(n794) );
  NOR2_X1 U410 ( .A1(n769), .A2(n220), .ZN(n1216) );
  NAND2_X1 U411 ( .A1(n216), .A2(n735), .ZN(n1198) );
  INV_X1 U412 ( .A(n676), .ZN(n1505) );
  AND2_X4 U413 ( .A1(n686), .A2(n684), .ZN(n462) );
  INV_X2 U414 ( .A(n526), .ZN(n503) );
  OR2_X4 U415 ( .A1(n395), .A2(n1551), .ZN(n790) );
  XOR2_X2 U416 ( .A(n739), .B(n740), .Z(n344) );
  XOR2_X1 U417 ( .A(n745), .B(n744), .Z(n346) );
  AOI21_X1 U418 ( .B1(n281), .B2(n646), .A(n644), .ZN(n714) );
  INV_X2 U419 ( .A(n1132), .ZN(n644) );
  OR2_X1 U420 ( .A1(n624), .A2(n623), .ZN(n401) );
  INV_X4 U423 ( .A(n688), .ZN(n400) );
  NOR2_X1 U424 ( .A1(n208), .A2(n247), .ZN(U6_Z_23) );
  NOR2_X1 U425 ( .A1(n208), .A2(n221), .ZN(U6_Z_24) );
  NOR2_X1 U426 ( .A1(n775), .A2(n823), .ZN(n1215) );
  INV_X4 U427 ( .A(in_b_mac[13]), .ZN(n442) );
  XNOR2_X1 U428 ( .A(n1489), .B(n1488), .ZN(n407) );
  XOR2_X1 U429 ( .A(n347), .B(n1501), .Z(n209) );
  XNOR2_X1 U430 ( .A(n286), .B(n1499), .ZN(n347) );
  XNOR2_X1 U431 ( .A(n1470), .B(n1474), .ZN(n279) );
  XOR2_X1 U432 ( .A(n1473), .B(n1472), .Z(n1474) );
  XNOR2_X1 U433 ( .A(n348), .B(n297), .ZN(n557) );
  XOR2_X1 U434 ( .A(n572), .B(n240), .Z(n348) );
  XOR2_X1 U435 ( .A(n349), .B(n1494), .Z(n217) );
  XNOR2_X1 U436 ( .A(n295), .B(n1492), .ZN(n349) );
  XNOR2_X1 U437 ( .A(n1497), .B(n350), .ZN(n212) );
  XOR2_X1 U438 ( .A(n1495), .B(n324), .Z(n350) );
  XNOR2_X1 U439 ( .A(n551), .B(n528), .ZN(n409) );
  XOR2_X1 U442 ( .A(n409), .B(n278), .Z(n534) );
  XOR2_X1 U443 ( .A(n351), .B(n530), .Z(n517) );
  XNOR2_X1 U444 ( .A(n262), .B(n234), .ZN(n351) );
  AND2_X4 U445 ( .A1(n246), .A2(U1_C_4_), .ZN(n547) );
  OAI21_X2 U446 ( .B1(U1_C_1_), .B2(n252), .A(n497), .ZN(n488) );
  AND2_X4 U447 ( .A1(n715), .A2(U1_C_8_), .ZN(n652) );
  INV_X4 U448 ( .A(in_a_mac[3]), .ZN(n1449) );
  XNOR2_X2 U449 ( .A(n353), .B(n1139), .ZN(n1125) );
  XNOR2_X2 U450 ( .A(n1135), .B(n1134), .ZN(n353) );
  NOR2_X2 U451 ( .A1(n1500), .A2(n1501), .ZN(n953) );
  XNOR2_X2 U452 ( .A(n354), .B(n1192), .ZN(n1487) );
  XNOR2_X2 U455 ( .A(n1193), .B(n1197), .ZN(n354) );
  XNOR2_X2 U456 ( .A(n355), .B(n1142), .ZN(n1476) );
  XNOR2_X2 U459 ( .A(n1143), .B(n1147), .ZN(n355) );
  XNOR2_X2 U461 ( .A(n356), .B(n1177), .ZN(n1484) );
  XNOR2_X2 U462 ( .A(n1179), .B(n1183), .ZN(n356) );
  XNOR2_X2 U463 ( .A(n357), .B(n1164), .ZN(n1479) );
  XNOR2_X2 U464 ( .A(n1163), .B(n1162), .ZN(n357) );
  XOR2_X2 U465 ( .A(n793), .B(n358), .Z(n1223) );
  XNOR2_X2 U466 ( .A(n1508), .B(n1530), .ZN(n358) );
  XNOR2_X2 U467 ( .A(n1206), .B(n359), .ZN(n1394) );
  XNOR2_X2 U468 ( .A(n389), .B(n1207), .ZN(n359) );
  XNOR2_X2 U469 ( .A(n363), .B(n1222), .ZN(n1398) );
  XNOR2_X2 U470 ( .A(n1223), .B(n1221), .ZN(n363) );
  XNOR2_X2 U471 ( .A(n1424), .B(n1423), .ZN(n1426) );
  OR2_X1 U472 ( .A1(n844), .A2(n364), .ZN(n1234) );
  AND2_X4 U473 ( .A1(n843), .A2(n1508), .ZN(n364) );
  AOI21_X2 U474 ( .B1(n845), .B2(n1530), .A(n793), .ZN(n844) );
  XOR2_X2 U475 ( .A(n365), .B(n313), .Z(n255) );
  XNOR2_X2 U476 ( .A(n1406), .B(n1405), .ZN(n365) );
  XNOR2_X2 U477 ( .A(n369), .B(n952), .ZN(n1498) );
  XNOR2_X2 U478 ( .A(n370), .B(n1127), .ZN(n1472) );
  XNOR2_X2 U479 ( .A(n1126), .B(n1125), .ZN(n370) );
  XNOR2_X2 U480 ( .A(n371), .B(n985), .ZN(n1138) );
  XNOR2_X2 U481 ( .A(n981), .B(n653), .ZN(n371) );
  XNOR2_X2 U482 ( .A(n372), .B(n679), .ZN(n705) );
  XNOR2_X2 U483 ( .A(n704), .B(n373), .ZN(n969) );
  XNOR2_X2 U484 ( .A(n703), .B(n702), .ZN(n373) );
  XNOR2_X2 U485 ( .A(n374), .B(n683), .ZN(n1040) );
  XNOR2_X2 U488 ( .A(n682), .B(n635), .ZN(n374) );
  XNOR2_X2 U489 ( .A(n376), .B(n673), .ZN(n1163) );
  XNOR2_X2 U490 ( .A(n672), .B(n1172), .ZN(n376) );
  XNOR2_X2 U491 ( .A(n377), .B(n1185), .ZN(n1179) );
  XNOR2_X2 U492 ( .A(n1186), .B(n343), .ZN(n377) );
  XNOR2_X2 U493 ( .A(n1155), .B(n378), .ZN(n1143) );
  XNOR2_X2 U494 ( .A(n1504), .B(n1503), .ZN(n378) );
  XNOR2_X2 U496 ( .A(n1463), .B(n379), .ZN(n1135) );
  XNOR2_X2 U497 ( .A(n656), .B(n657), .ZN(n379) );
  AOI21_X1 U498 ( .B1(n754), .B2(n751), .A(n1538), .ZN(n808) );
  XNOR2_X2 U499 ( .A(n733), .B(n381), .ZN(n1193) );
  XNOR2_X2 U500 ( .A(n735), .B(n216), .ZN(n381) );
  XNOR2_X2 U501 ( .A(n382), .B(n456), .ZN(n698) );
  XNOR2_X2 U502 ( .A(n455), .B(n783), .ZN(n382) );
  XNOR2_X2 U503 ( .A(n383), .B(n384), .ZN(n701) );
  XNOR2_X2 U504 ( .A(n1462), .B(n779), .ZN(n384) );
  AND2_X1 U505 ( .A1(n474), .A2(n653), .ZN(n473) );
  AND2_X1 U506 ( .A1(n779), .A2(n777), .ZN(n1456) );
  AND2_X1 U507 ( .A1(n864), .A2(n862), .ZN(n1448) );
  XOR2_X2 U508 ( .A(n840), .B(n386), .Z(n1237) );
  XOR2_X2 U509 ( .A(n841), .B(n842), .Z(n386) );
  AOI21_X1 U510 ( .B1(n731), .B2(n732), .A(n1506), .ZN(n769) );
  AOI21_X2 U511 ( .B1(n1509), .B2(n848), .A(n889), .ZN(n841) );
  AOI21_X2 U512 ( .B1(n890), .B2(n1527), .A(n847), .ZN(n889) );
  XOR2_X2 U513 ( .A(n862), .B(n387), .Z(n795) );
  XNOR2_X2 U514 ( .A(n1453), .B(n864), .ZN(n387) );
  AOI21_X2 U515 ( .B1(n911), .B2(n908), .A(n1536), .ZN(n887) );
  OAI21_X2 U516 ( .B1(n908), .B2(n911), .A(n910), .ZN(n941) );
  AOI21_X1 U517 ( .B1(n803), .B2(n800), .A(n1545), .ZN(n797) );
  OAI21_X1 U518 ( .B1(n800), .B2(n803), .A(n802), .ZN(n870) );
  AOI21_X1 U519 ( .B1(n805), .B2(n806), .A(n1531), .ZN(n798) );
  XOR2_X2 U520 ( .A(n1439), .B(n1438), .Z(n388) );
  OAI21_X1 U521 ( .B1(n216), .B2(n735), .A(n733), .ZN(n770) );
  OAI21_X1 U522 ( .B1(n765), .B2(n764), .A(n762), .ZN(n849) );
  OAI21_X1 U523 ( .B1(n1505), .B2(n707), .A(n674), .ZN(n706) );
  XNOR2_X2 U524 ( .A(n766), .B(n390), .ZN(n389) );
  XNOR2_X2 U525 ( .A(n220), .B(n769), .ZN(n390) );
  AOI21_X2 U526 ( .B1(n973), .B2(n970), .A(n1535), .ZN(n920) );
  OAI21_X2 U527 ( .B1(n970), .B2(n973), .A(n972), .ZN(n1008) );
  AOI21_X2 U528 ( .B1(n1000), .B2(n997), .A(n1534), .ZN(n988) );
  OAI21_X2 U529 ( .B1(n997), .B2(n1000), .A(n999), .ZN(n1057) );
  OAI21_X2 U532 ( .B1(n924), .B2(n1515), .A(n922), .ZN(n962) );
  OAI21_X2 U533 ( .B1(n1540), .B2(n1032), .A(n1063), .ZN(n1026) );
  OAI21_X2 U537 ( .B1(n1031), .B2(n1526), .A(n1033), .ZN(n1063) );
  OAI21_X2 U538 ( .B1(n996), .B2(n1518), .A(n958), .ZN(n995) );
  OAI21_X2 U539 ( .B1(n1085), .B2(n1539), .A(n1100), .ZN(n1077) );
  OAI21_X2 U540 ( .B1(n1101), .B2(n1525), .A(n1086), .ZN(n1100) );
  XNOR2_X2 U541 ( .A(n882), .B(n901), .ZN(n391) );
  XNOR2_X2 U543 ( .A(n713), .B(n392), .ZN(n743) );
  XNOR2_X2 U544 ( .A(n712), .B(n711), .ZN(n392) );
  XNOR2_X2 U545 ( .A(n393), .B(n568), .ZN(n573) );
  XNOR2_X2 U547 ( .A(n394), .B(n342), .ZN(n703) );
  XNOR2_X2 U548 ( .A(n1017), .B(n1040), .ZN(n394) );
  OAI21_X2 U549 ( .B1(n533), .B2(n532), .A(n531), .ZN(n550) );
  NOR2_X2 U550 ( .A1(n1383), .A2(n1382), .ZN(n1385) );
  XNOR2_X2 U551 ( .A(n1384), .B(n1381), .ZN(n396) );
  XNOR2_X2 U552 ( .A(n397), .B(n1166), .ZN(n676) );
  XNOR2_X2 U553 ( .A(n1167), .B(n1168), .ZN(n397) );
  XOR2_X2 U554 ( .A(n398), .B(n1014), .Z(n697) );
  XNOR2_X2 U558 ( .A(n987), .B(n1004), .ZN(n398) );
  XNOR2_X2 U559 ( .A(n399), .B(n621), .ZN(n1126) );
  XNOR2_X2 U560 ( .A(n624), .B(n623), .ZN(n399) );
  NAND2_X2 U561 ( .A1(n400), .A2(n401), .ZN(n1153) );
  AND2_X1 U566 ( .A1(n694), .A2(n745), .ZN(n693) );
  XNOR2_X2 U567 ( .A(n1379), .B(n1378), .ZN(n1366) );
  AOI21_X2 U568 ( .B1(n879), .B2(n878), .A(n876), .ZN(n967) );
  AOI21_X2 U569 ( .B1(n1511), .B2(n1517), .A(n791), .ZN(n907) );
  AOI21_X2 U570 ( .B1(n868), .B2(n360), .A(n1554), .ZN(n806) );
  OAI21_X1 U572 ( .B1(n808), .B2(n739), .A(n809), .ZN(n731) );
  OAI21_X1 U574 ( .B1(n1507), .B2(n1537), .A(n740), .ZN(n809) );
  AOI21_X2 U575 ( .B1(n854), .B2(n1514), .A(n1510), .ZN(n890) );
  OAI21_X2 U576 ( .B1(n1514), .B2(n854), .A(n423), .ZN(n895) );
  XOR2_X2 U577 ( .A(n403), .B(n698), .Z(n1178) );
  XNOR2_X2 U578 ( .A(n1173), .B(n701), .ZN(n403) );
  AOI21_X2 U579 ( .B1(n837), .B2(n835), .A(n1516), .ZN(n883) );
  OAI21_X2 U580 ( .B1(n835), .B2(n837), .A(n838), .ZN(n930) );
  XNOR2_X2 U581 ( .A(n774), .B(n775), .ZN(n404) );
  AOI21_X1 U582 ( .B1(n823), .B2(n775), .A(n774), .ZN(n822) );
  OR2_X1 U583 ( .A1(n405), .A2(n896), .ZN(n606) );
  AND2_X4 U585 ( .A1(n716), .A2(n717), .ZN(n405) );
  INV_X4 U586 ( .A(in_b_mac[14]), .ZN(n441) );
  OAI21_X2 U587 ( .B1(n1542), .B2(n899), .A(n946), .ZN(n885) );
  OAI21_X2 U588 ( .B1(n1513), .B2(n947), .A(n913), .ZN(n946) );
  AOI21_X2 U591 ( .B1(n885), .B2(n1256), .A(n940), .ZN(n1502) );
  AOI21_X2 U592 ( .B1(n1512), .B2(n888), .A(n887), .ZN(n940) );
  OAI21_X2 U593 ( .B1(n964), .B2(n965), .A(n966), .ZN(n1012) );
  OAI21_X2 U594 ( .B1(n926), .B2(n929), .A(n928), .ZN(n978) );
  AOI21_X2 U597 ( .B1(n957), .B2(n956), .A(n954), .ZN(n1034) );
  OR2_X1 U598 ( .A1(n406), .A2(n1056), .ZN(n1526) );
  AND2_X4 U599 ( .A1(n430), .A2(n1442), .ZN(n406) );
  OAI21_X2 U600 ( .B1(n1529), .B2(n988), .A(n1521), .ZN(n1027) );
  AOI21_X2 U601 ( .B1(n988), .B2(n1529), .A(n990), .ZN(n1053) );
  OAI21_X2 U602 ( .B1(n994), .B2(n993), .A(n991), .ZN(n1028) );
  OAI21_X2 U605 ( .B1(n1027), .B2(n1026), .A(n1024), .ZN(n1049) );
  OAI21_X2 U606 ( .B1(n1021), .B2(n1022), .A(n1023), .ZN(n1067) );
  XOR2_X2 U607 ( .A(n407), .B(n429), .Z(n259) );
  AOI21_X2 U608 ( .B1(n1048), .B2(n1047), .A(n1045), .ZN(n1081) );
  AOI21_X1 U609 ( .B1(n721), .B2(n438), .A(n1111), .ZN(n1095) );
  AOI21_X2 U610 ( .B1(n1094), .B2(n1532), .A(n1095), .ZN(n1110) );
  OAI21_X2 U611 ( .B1(n1077), .B2(n1080), .A(n1079), .ZN(n1097) );
  OR2_X1 U614 ( .A1(n408), .A2(n1123), .ZN(n634) );
  AND2_X4 U615 ( .A1(n814), .A2(n437), .ZN(n408) );
  AND2_X1 U617 ( .A1(n828), .A2(U1_C_6_), .ZN(n827) );
  XNOR2_X2 U618 ( .A(n410), .B(n681), .ZN(n1017) );
  XNOR2_X2 U622 ( .A(n680), .B(U1_C_10_), .ZN(n410) );
  XNOR2_X2 U623 ( .A(n411), .B(n385), .ZN(n772) );
  XNOR2_X2 U624 ( .A(n412), .B(n402), .ZN(n865) );
  XNOR2_X2 U625 ( .A(n715), .B(U1_C_8_), .ZN(n412) );
  XNOR2_X2 U626 ( .A(n287), .B(U1_C_4_), .ZN(n413) );
  XNOR2_X2 U628 ( .A(n513), .B(U1_C_2_), .ZN(n414) );
  INV_X4 U629 ( .A(in_a_mac[9]), .ZN(n435) );
  XNOR2_X2 U632 ( .A(n1449), .B(in_a_mac[4]), .ZN(n418) );
  XNOR2_X2 U633 ( .A(n420), .B(n483), .ZN(n1132) );
  XNOR2_X2 U634 ( .A(n482), .B(U1_C_12_), .ZN(n420) );
  OAI21_X2 U635 ( .B1(U1_C_11_), .B2(n484), .A(n1129), .ZN(n621) );
  XNOR2_X2 U640 ( .A(in_a_mac[12]), .B(n1552), .ZN(n421) );
  XNOR2_X2 U641 ( .A(n422), .B(n618), .ZN(n1173) );
  XNOR2_X2 U642 ( .A(n615), .B(U1_C_14_), .ZN(n422) );
  INV_X4 U643 ( .A(in_a_mac[13]), .ZN(n1553) );
  INV_X4 U644 ( .A(in_a_mac[15]), .ZN(n1554) );
  AOI21_X2 U645 ( .B1(n898), .B2(U1_C_16_), .A(n899), .ZN(n897) );
  AND2_X1 U646 ( .A1(U1_C_15_), .A2(n1444), .ZN(n423) );
  OAI21_X2 U647 ( .B1(n1541), .B2(n65), .A(n979), .ZN(n928) );
  OAI21_X2 U649 ( .B1(U1_C_17_), .B2(n932), .A(U1_C_18_), .ZN(n979) );
  AOI21_X2 U650 ( .B1(n1007), .B2(n593), .A(n1519), .ZN(n957) );
  OAI21_X2 U651 ( .B1(n593), .B2(n1007), .A(U1_C_20_), .ZN(n1038) );
  AOI21_X2 U652 ( .B1(n1037), .B2(n1035), .A(n1522), .ZN(n990) );
  OAI21_X2 U655 ( .B1(n1035), .B2(n1037), .A(n41), .ZN(n1054) );
  AOI21_X2 U656 ( .B1(n1052), .B2(n1050), .A(n1523), .ZN(n1047) );
  OAI21_X2 U657 ( .B1(n1050), .B2(n1052), .A(n29), .ZN(n1087) );
  OAI21_X2 U658 ( .B1(n1533), .B2(n41), .A(n1069), .ZN(n1021) );
  OAI21_X2 U659 ( .B1(U1_C_21_), .B2(n1070), .A(U1_C_22_), .ZN(n1069) );
  OAI21_X2 U664 ( .B1(n1528), .B2(n29), .A(n1098), .ZN(n1079) );
  OAI21_X2 U665 ( .B1(U1_C_23_), .B2(n1083), .A(U1_C_24_), .ZN(n1098) );
  AOI21_X2 U666 ( .B1(n1076), .B2(n1074), .A(n1524), .ZN(n1094) );
  OAI21_X2 U667 ( .B1(n1074), .B2(n1076), .A(n18), .ZN(n1112) );
  OAI21_X2 U668 ( .B1(U1_C_25_), .B2(n1092), .A(U1_C_26_), .ZN(n1116) );
  OAI21_X2 U670 ( .B1(U1_C_27_), .B2(n367), .A(U1_C_28_), .ZN(n366) );
  OAI21_X2 U672 ( .B1(n1107), .B2(n1109), .A(n12), .ZN(n1121) );
  INV_X4 U673 ( .A(n485), .ZN(n208) );
  NAND2_X2 U675 ( .A1(n834), .A2(n832), .ZN(n839) );
  NOR2_X2 U676 ( .A1(n1420), .A2(n1297), .ZN(n1302) );
  OAI22_X2 U679 ( .A1(n1291), .A2(n1417), .B1(n1290), .B2(n1415), .ZN(n1420)
         );
  OAI22_X1 U680 ( .A1(n236), .A2(n626), .B1(n625), .B2(n268), .ZN(n629) );
  AOI21_X1 U682 ( .B1(n236), .B2(n268), .A(n626), .ZN(n1443) );
  OAI22_X1 U683 ( .A1(n236), .A2(n625), .B1(n1450), .B2(n268), .ZN(n1199) );
  OAI22_X1 U684 ( .A1(n236), .A2(n1450), .B1(n1455), .B2(n268), .ZN(n1461) );
  OAI22_X1 U685 ( .A1(n236), .A2(n1455), .B1(n1454), .B2(n268), .ZN(n1462) );
  OAI22_X1 U686 ( .A1(n1148), .A2(n268), .B1(n236), .B2(n1454), .ZN(n1457) );
  OAI22_X1 U691 ( .A1(n236), .A2(n1148), .B1(n977), .B2(n268), .ZN(n1151) );
  OAI22_X1 U692 ( .A1(n236), .A2(n977), .B1(n974), .B2(n268), .ZN(n1463) );
  OAI22_X1 U693 ( .A1(n236), .A2(n974), .B1(n662), .B2(n253), .ZN(n481) );
  INV_X1 U697 ( .A(n432), .ZN(n502) );
  NOR2_X1 U700 ( .A1(n768), .A2(n767), .ZN(n771) );
  AOI21_X1 U702 ( .B1(n280), .B2(n440), .A(n1089), .ZN(n1085) );
  OAI22_X1 U703 ( .A1(n440), .A2(n1089), .B1(n1062), .B2(n280), .ZN(n1052) );
  OAI22_X1 U704 ( .A1(n440), .A2(n1062), .B1(n1055), .B2(n280), .ZN(n1061) );
  OAI22_X1 U705 ( .A1(n440), .A2(n1055), .B1(n1039), .B2(n280), .ZN(n1035) );
  OAI22_X1 U706 ( .A1(n440), .A2(n1039), .B1(n1011), .B2(n280), .ZN(n1007) );
  OAI22_X1 U707 ( .A1(n440), .A2(n980), .B1(n949), .B2(n280), .ZN(n932) );
  OAI22_X1 U708 ( .A1(n440), .A2(n1011), .B1(n980), .B2(n280), .ZN(n973) );
  OAI22_X1 U709 ( .A1(n440), .A2(n949), .B1(n900), .B2(n280), .ZN(n947) );
  OAI22_X1 U710 ( .A1(n440), .A2(n900), .B1(n873), .B2(n280), .ZN(n854) );
  OAI22_X1 U711 ( .A1(n440), .A2(n873), .B1(n829), .B2(n280), .ZN(n800) );
  OAI22_X1 U712 ( .A1(n440), .A2(n829), .B1(n816), .B2(n280), .ZN(n783) );
  OAI22_X1 U714 ( .A1(n440), .A2(n816), .B1(n757), .B2(n280), .ZN(n811) );
  OAI22_X1 U715 ( .A1(n440), .A2(n757), .B1(n722), .B2(n280), .ZN(n684) );
  OAI22_X1 U716 ( .A1(n640), .A2(n440), .B1(n280), .B2(n689), .ZN(n694) );
  OAI22_X1 U718 ( .A1(n950), .A2(n952), .B1(n749), .B2(n938), .ZN(n968) );
  INV_X4 U719 ( .A(n635), .ZN(n425) );
  XOR2_X1 U720 ( .A(n1437), .B(n228), .Z(n243) );
  OAI22_X2 U721 ( .A1(n1411), .A2(n1279), .B1(n1278), .B2(n1277), .ZN(n1416)
         );
  OAI22_X1 U724 ( .A1(n713), .A2(n667), .B1(n270), .B2(n666), .ZN(n704) );
  XNOR2_X1 U725 ( .A(n1433), .B(n311), .ZN(n244) );
  XNOR2_X1 U728 ( .A(n1410), .B(n328), .ZN(n250) );
  NOR2_X1 U730 ( .A1(n415), .A2(n221), .ZN(U5_Z_8) );
  NOR2_X1 U731 ( .A1(n415), .A2(n242), .ZN(U5_Z_12) );
  NOR2_X1 U732 ( .A1(n415), .A2(n244), .ZN(U5_Z_10) );
  NOR2_X1 U733 ( .A1(n415), .A2(n245), .ZN(U5_Z_9) );
  NOR2_X1 U734 ( .A1(n415), .A2(n250), .ZN(U5_Z_4) );
  NOR2_X1 U735 ( .A1(n247), .A2(n415), .ZN(U5_Z_7) );
  NOR2_X1 U736 ( .A1(n248), .A2(n415), .ZN(U5_Z_6) );
  NOR2_X1 U738 ( .A1(n257), .A2(n415), .ZN(U5_Z_1) );
  NOR2_X1 U739 ( .A1(n415), .A2(n255), .ZN(U5_Z_3) );
  NOR2_X1 U742 ( .A1(n243), .A2(n415), .ZN(U5_Z_11) );
  NOR2_X1 U744 ( .A1(n249), .A2(n415), .ZN(U5_Z_5) );
  NOR2_X1 U745 ( .A1(n256), .A2(n415), .ZN(U5_Z_2) );
  NOR2_X1 U746 ( .A1(n258), .A2(n415), .ZN(U5_Z_0) );
  NAND2_X1 U747 ( .A1(n431), .A2(n273), .ZN(n583) );
  OAI22_X1 U748 ( .A1(n627), .A2(n273), .B1(n431), .B2(n602), .ZN(n605) );
  OAI22_X1 U751 ( .A1(n431), .A2(n588), .B1(n602), .B2(n273), .ZN(n589) );
  OAI22_X1 U752 ( .A1(n431), .A2(n1446), .B1(n450), .B2(n273), .ZN(n447) );
  OAI22_X1 U753 ( .A1(n431), .A2(n627), .B1(n1447), .B2(n273), .ZN(n1211) );
  OAI22_X1 U755 ( .A1(n431), .A2(n1447), .B1(n1446), .B2(n273), .ZN(n1453) );
  OAI22_X1 U757 ( .A1(n431), .A2(n450), .B1(n470), .B2(n273), .ZN(n453) );
  OAI22_X1 U758 ( .A1(n471), .A2(n273), .B1(n431), .B2(n470), .ZN(n1166) );
  OAI22_X1 U762 ( .A1(n431), .A2(n471), .B1(n472), .B2(n273), .ZN(n459) );
  OAI22_X1 U763 ( .A1(n431), .A2(n472), .B1(n669), .B2(n273), .ZN(n474) );
  OAI22_X1 U766 ( .A1(n431), .A2(n669), .B1(n687), .B2(n273), .ZN(n987) );
  OAI22_X1 U767 ( .A1(n431), .A2(n687), .B1(n685), .B2(n1445), .ZN(n745) );
  OAI22_X1 U772 ( .A1(n431), .A2(n727), .B1(n723), .B2(n1445), .ZN(n788) );
  OAI22_X1 U774 ( .A1(n431), .A2(n685), .B1(n727), .B2(n1445), .ZN(n658) );
  NAND2_X1 U775 ( .A1(n543), .A2(n1445), .ZN(n544) );
  XOR2_X1 U778 ( .A(n263), .B(n1466), .Z(n1468) );
  INV_X4 U779 ( .A(n784), .ZN(n426) );
  NOR2_X1 U780 ( .A1(n260), .A2(n742), .ZN(n749) );
  XNOR2_X1 U782 ( .A(n1478), .B(n276), .ZN(n274) );
  INV_X1 U783 ( .A(n266), .ZN(n528) );
  OAI22_X1 U786 ( .A1(n540), .A2(n539), .B1(n537), .B2(n538), .ZN(n572) );
  INV_X1 U787 ( .A(n1471), .ZN(n1473) );
  INV_X1 U788 ( .A(n1420), .ZN(n1303) );
  INV_X2 U790 ( .A(n1449), .ZN(n428) );
  NOR2_X1 U792 ( .A1(n415), .A2(n215), .ZN(U5_Z_13) );
  XOR2_X1 U793 ( .A(n1396), .B(n336), .Z(n258) );
  XNOR2_X1 U798 ( .A(n1404), .B(n1403), .ZN(n256) );
  XOR2_X1 U799 ( .A(in_a_mac[7]), .B(in_a_mac[6]), .Z(n1066) );
  XOR2_X1 U802 ( .A(n299), .B(n1481), .Z(n269) );
  XNOR2_X1 U803 ( .A(n1486), .B(n337), .ZN(n264) );
  XNOR2_X1 U804 ( .A(n1398), .B(n291), .ZN(n1400) );
  XOR2_X1 U806 ( .A(n290), .B(n1427), .Z(n1430) );
  XOR2_X1 U807 ( .A(n288), .B(n1419), .Z(n1422) );
  XOR2_X1 U808 ( .A(n289), .B(n1415), .Z(n1418) );
  XOR2_X1 U812 ( .A(n755), .B(n759), .Z(n580) );
  OAI22_X1 U813 ( .A1(n787), .A2(n786), .B1(n785), .B2(n784), .ZN(n856) );
  NAND2_X4 U814 ( .A1(n1066), .A2(n430), .ZN(n1442) );
  INV_X4 U815 ( .A(n446), .ZN(n463) );
  INV_X4 U816 ( .A(n447), .ZN(n465) );
  NOR2_X2 U817 ( .A1(n447), .A2(n446), .ZN(n449) );
  XOR2_X2 U818 ( .A(n1444), .B(U1_C_15_), .Z(n464) );
  INV_X4 U820 ( .A(n464), .ZN(n448) );
  OAI22_X2 U821 ( .A1(n463), .A2(n465), .B1(n449), .B2(n448), .ZN(n764) );
  INV_X4 U824 ( .A(n453), .ZN(n456) );
  INV_X4 U825 ( .A(n783), .ZN(n451) );
  NOR2_X2 U826 ( .A1(n456), .A2(n451), .ZN(n452) );
  OAI22_X2 U827 ( .A1(n783), .A2(n453), .B1(n452), .B2(n455), .ZN(n823) );
  INV_X4 U828 ( .A(n361), .ZN(n454) );
  INV_X4 U830 ( .A(n622), .ZN(n618) );
  INV_X4 U832 ( .A(n1173), .ZN(n700) );
  NOR2_X2 U833 ( .A1(n698), .A2(n700), .ZN(n457) );
  OR2_X1 U840 ( .A1(n776), .A2(n457), .ZN(n735) );
  OAI22_X2 U842 ( .A1(n747), .A2(n717), .B1(n696), .B2(n716), .ZN(n484) );
  NAND2_X2 U843 ( .A1(U1_C_11_), .A2(n484), .ZN(n1129) );
  INV_X4 U848 ( .A(n1129), .ZN(n460) );
  INV_X4 U850 ( .A(n459), .ZN(n1130) );
  NOR2_X2 U851 ( .A1(n1130), .A2(n1129), .ZN(n458) );
  OAI22_X2 U852 ( .A1(n460), .A2(n459), .B1(n458), .B2(n1128), .ZN(n672) );
  XOR2_X2 U853 ( .A(n352), .B(in_b_mac[10]), .Z(n1148) );
  XOR2_X2 U854 ( .A(n352), .B(in_b_mac[9]), .Z(n977) );
  OAI22_X2 U857 ( .A1(n684), .A2(n686), .B1(n462), .B2(n1151), .ZN(n673) );
  XOR2_X2 U858 ( .A(n464), .B(n463), .Z(n466) );
  XOR2_X2 U863 ( .A(n466), .B(n465), .Z(n733) );
  OAI22_X2 U864 ( .A1(n817), .A2(n717), .B1(n746), .B2(n716), .ZN(n1460) );
  XOR2_X2 U865 ( .A(n1460), .B(U1_C_13_), .Z(n1167) );
  INV_X4 U867 ( .A(n468), .ZN(n483) );
  NOR2_X2 U869 ( .A1(n468), .A2(n467), .ZN(n469) );
  OAI22_X2 U870 ( .A1(n746), .A2(n717), .B1(n747), .B2(n716), .ZN(n482) );
  OAI22_X2 U875 ( .A1(U1_C_12_), .A2(n483), .B1(n469), .B2(n482), .ZN(n1168)
         );
  INV_X4 U876 ( .A(n1166), .ZN(n1171) );
  INV_X4 U879 ( .A(n474), .ZN(n985) );
  OAI22_X2 U881 ( .A1(n653), .A2(n474), .B1(n473), .B2(n981), .ZN(n646) );
  NOR2_X2 U882 ( .A1(n281), .A2(n646), .ZN(n475) );
  OR2_X1 U883 ( .A1(n714), .A2(n475), .ZN(n707) );
  OAI22_X2 U885 ( .A1(n696), .A2(n717), .B1(n660), .B2(n716), .ZN(n479) );
  INV_X4 U887 ( .A(n680), .ZN(n478) );
  INV_X4 U888 ( .A(n479), .ZN(n681) );
  NOR2_X2 U889 ( .A1(n681), .A2(n476), .ZN(n477) );
  OAI22_X2 U890 ( .A1(U1_C_10_), .A2(n479), .B1(n478), .B2(n477), .ZN(n623) );
  XOR2_X2 U893 ( .A(n352), .B(in_b_mac[8]), .Z(n974) );
  XOR2_X2 U894 ( .A(n427), .B(in_b_mac[7]), .Z(n662) );
  INV_X4 U899 ( .A(n481), .ZN(n683) );
  NOR2_X2 U901 ( .A1(n683), .A2(n425), .ZN(n480) );
  OAI22_X2 U903 ( .A1(n692), .A2(n430), .B1(n665), .B2(n1442), .ZN(n682) );
  OAI22_X2 U906 ( .A1(n635), .A2(n481), .B1(n480), .B2(n682), .ZN(n624) );
  OR4_X1 U907 ( .A1(bitselect1[1]), .A2(bitselect1[0]), .A3(bitselect1[3]), 
        .A4(bitselect1[2]), .ZN(n485) );
  XOR2_X2 U908 ( .A(n491), .B(U1_C_0_), .Z(n486) );
  NOR2_X2 U910 ( .A1(n208), .A2(n486), .ZN(U6_Z_0) );
  NAND2_X2 U911 ( .A1(n487), .A2(U1_C_1_), .ZN(n497) );
  INV_X4 U912 ( .A(n488), .ZN(n493) );
  NOR2_X2 U913 ( .A1(n318), .A2(n444), .ZN(n489) );
  NAND2_X2 U914 ( .A1(n493), .A2(n492), .ZN(n498) );
  NOR3_X2 U918 ( .A1(n495), .A2(n494), .A3(n208), .ZN(U6_Z_1) );
  XOR2_X2 U922 ( .A(n433), .B(in_b_mac[2]), .Z(n506) );
  OAI22_X2 U925 ( .A1(n506), .A2(n717), .B1(n496), .B2(n716), .ZN(n516) );
  INV_X4 U926 ( .A(n516), .ZN(n513) );
  NAND2_X2 U929 ( .A1(n498), .A2(n497), .ZN(n509) );
  XNOR2_X2 U930 ( .A(n510), .B(n509), .ZN(n499) );
  NOR2_X2 U931 ( .A1(n208), .A2(n499), .ZN(U6_Z_2) );
  NAND2_X2 U935 ( .A1(n502), .A2(n444), .ZN(n500) );
  NAND2_X2 U936 ( .A1(n500), .A2(n254), .ZN(n501) );
  NAND2_X2 U938 ( .A1(n428), .A2(n501), .ZN(n519) );
  XOR2_X2 U945 ( .A(n427), .B(in_b_mac[1]), .Z(n526) );
  NAND2_X2 U947 ( .A1(n503), .A2(n502), .ZN(n504) );
  XNOR2_X2 U949 ( .A(n523), .B(n519), .ZN(n508) );
  NAND2_X2 U950 ( .A1(n507), .A2(U1_C_3_), .ZN(n535) );
  XNOR2_X2 U951 ( .A(n508), .B(n518), .ZN(n532) );
  NAND2_X2 U952 ( .A1(n510), .A2(n509), .ZN(n529) );
  INV_X4 U953 ( .A(n511), .ZN(n515) );
  NOR2_X2 U954 ( .A1(n513), .A2(n512), .ZN(n514) );
  NOR2_X2 U955 ( .A1(n208), .A2(n517), .ZN(U6_Z_3) );
  INV_X4 U956 ( .A(n519), .ZN(n524) );
  INV_X4 U957 ( .A(n518), .ZN(n522) );
  NOR2_X2 U958 ( .A1(n520), .A2(n519), .ZN(n521) );
  OAI22_X2 U959 ( .A1(n524), .A2(n271), .B1(n522), .B2(n521), .ZN(n551) );
  XOR2_X2 U960 ( .A(n352), .B(in_b_mac[2]), .Z(n545) );
  INV_X4 U961 ( .A(n539), .ZN(n536) );
  XNOR2_X2 U962 ( .A(n527), .B(n536), .ZN(n552) );
  NOR2_X2 U963 ( .A1(n529), .A2(n530), .ZN(n533) );
  NAND2_X2 U964 ( .A1(n529), .A2(n530), .ZN(n531) );
  NOR2_X2 U965 ( .A1(n208), .A2(n534), .ZN(U6_Z_4) );
  NOR2_X2 U966 ( .A1(n536), .A2(n535), .ZN(n537) );
  OAI22_X2 U967 ( .A1(n236), .A2(n565), .B1(n545), .B2(n254), .ZN(n558) );
  INV_X4 U968 ( .A(n551), .ZN(n549) );
  NAND2_X2 U969 ( .A1(n548), .A2(n549), .ZN(n556) );
  NAND2_X2 U970 ( .A1(n550), .A2(n551), .ZN(n554) );
  NAND2_X2 U971 ( .A1(n553), .A2(n554), .ZN(n555) );
  NOR2_X2 U972 ( .A1(n208), .A2(n557), .ZN(U6_Z_5) );
  OAI22_X2 U973 ( .A1(n574), .A2(n717), .B1(n559), .B2(n716), .ZN(n828) );
  INV_X4 U974 ( .A(n430), .ZN(n718) );
  OAI22_X2 U975 ( .A1(n431), .A2(n723), .B1(n564), .B2(n1445), .ZN(n784) );
  OAI22_X2 U976 ( .A1(n236), .A2(n819), .B1(n565), .B2(n253), .ZN(n786) );
  INV_X4 U977 ( .A(n786), .ZN(n782) );
  INV_X4 U978 ( .A(n767), .ZN(n778) );
  INV_X4 U979 ( .A(n568), .ZN(n570) );
  INV_X4 U980 ( .A(n752), .ZN(n759) );
  INV_X4 U981 ( .A(n572), .ZN(n576) );
  INV_X4 U982 ( .A(n573), .ZN(n575) );
  NOR2_X2 U983 ( .A1(n208), .A2(n581), .ZN(U6_Z_6) );
  INV_X4 U984 ( .A(n1526), .ZN(n1032) );
  INV_X4 U985 ( .A(n588), .ZN(n582) );
  NAND2_X2 U986 ( .A1(n583), .A2(n582), .ZN(n586) );
  INV_X4 U987 ( .A(n586), .ZN(n1260) );
  INV_X4 U988 ( .A(n1003), .ZN(n584) );
  NOR2_X2 U989 ( .A1(n1260), .A2(n584), .ZN(n585) );
  OAI22_X2 U990 ( .A1(n1003), .A2(n586), .B1(n585), .B2(n1259), .ZN(n956) );
  NOR2_X2 U991 ( .A1(n957), .A2(n956), .ZN(n587) );
  OR2_X1 U992 ( .A1(n1034), .A2(n587), .ZN(n993) );
  INV_X4 U993 ( .A(n589), .ZN(n600) );
  INV_X4 U994 ( .A(n599), .ZN(n592) );
  NOR2_X2 U995 ( .A1(n52), .A2(n589), .ZN(n591) );
  OAI22_X2 U996 ( .A1(n600), .A2(n593), .B1(n592), .B2(n591), .ZN(n964) );
  NAND2_X2 U997 ( .A1(n965), .A2(n964), .ZN(n594) );
  NAND2_X2 U998 ( .A1(n1012), .A2(n594), .ZN(n1518) );
  INV_X4 U999 ( .A(n939), .ZN(n598) );
  XOR2_X2 U1000 ( .A(n352), .B(in_b_mac[15]), .Z(n626) );
  NOR2_X2 U1001 ( .A1(n939), .A2(n982), .ZN(n597) );
  OAI22_X2 U1002 ( .A1(n598), .A2(n1544), .B1(n1443), .B2(n597), .ZN(n926) );
  XOR2_X2 U1003 ( .A(n599), .B(n593), .Z(n601) );
  XOR2_X2 U1004 ( .A(n601), .B(n600), .Z(n1240) );
  INV_X4 U1005 ( .A(n1240), .ZN(n876) );
  INV_X4 U1006 ( .A(n605), .ZN(n611) );
  INV_X4 U1007 ( .A(n935), .ZN(n603) );
  NOR2_X2 U1008 ( .A1(n611), .A2(n603), .ZN(n604) );
  OAI22_X2 U1009 ( .A1(n935), .A2(n605), .B1(n604), .B2(n610), .ZN(n878) );
  INV_X4 U1010 ( .A(n606), .ZN(n1200) );
  XOR2_X2 U1011 ( .A(n352), .B(in_b_mac[14]), .Z(n625) );
  XOR2_X2 U1012 ( .A(n427), .B(in_b_mac[13]), .Z(n1450) );
  INV_X4 U1013 ( .A(n1199), .ZN(n608) );
  NOR2_X2 U1014 ( .A1(n903), .A2(n606), .ZN(n607) );
  OAI22_X2 U1015 ( .A1(n1546), .A2(n1200), .B1(n608), .B2(n607), .ZN(n848) );
  NAND2_X2 U1016 ( .A1(n765), .A2(n764), .ZN(n609) );
  NAND2_X2 U1017 ( .A1(n849), .A2(n609), .ZN(n1508) );
  XOR2_X2 U1018 ( .A(n610), .B(n935), .Z(n612) );
  XOR2_X2 U1019 ( .A(n612), .B(n611), .Z(n1229) );
  INV_X4 U1020 ( .A(n1229), .ZN(n835) );
  INV_X4 U1021 ( .A(n615), .ZN(n620) );
  NOR2_X2 U1022 ( .A1(n618), .A2(n617), .ZN(n619) );
  OAI22_X2 U1023 ( .A1(U1_C_14_), .A2(n622), .B1(n620), .B2(n619), .ZN(n775)
         );
  INV_X4 U1024 ( .A(n629), .ZN(n1212) );
  NOR2_X2 U1025 ( .A1(n1212), .A2(U1_C_17_), .ZN(n628) );
  OAI22_X2 U1026 ( .A1(n65), .A2(n629), .B1(n628), .B2(n1211), .ZN(n888) );
  NAND2_X2 U1027 ( .A1(n929), .A2(n926), .ZN(n630) );
  NAND2_X2 U1028 ( .A1(n978), .A2(n630), .ZN(n1515) );
  NOR2_X2 U1029 ( .A1(n879), .A2(n878), .ZN(n631) );
  OR2_X1 U1030 ( .A1(n967), .A2(n631), .ZN(n924) );
  INV_X4 U1031 ( .A(n634), .ZN(n1361) );
  INV_X4 U1032 ( .A(n367), .ZN(n632) );
  XOR2_X2 U1033 ( .A(n632), .B(n1119), .Z(n1360) );
  INV_X4 U1034 ( .A(n1360), .ZN(n637) );
  NAND2_X2 U1035 ( .A1(n1109), .A2(n1107), .ZN(n633) );
  NOR2_X2 U1036 ( .A1(n1360), .A2(n634), .ZN(n636) );
  OAI22_X2 U1037 ( .A1(n1361), .A2(n637), .B1(n224), .B2(n636), .ZN(n1379) );
  OAI22_X2 U1038 ( .A1(n368), .A2(n360), .B1(n362), .B2(n361), .ZN(n1371) );
  NAND2_X2 U1039 ( .A1(n367), .A2(U1_C_27_), .ZN(n638) );
  NAND2_X2 U1040 ( .A1(n366), .A2(n638), .ZN(n1369) );
  INV_X4 U1041 ( .A(n1369), .ZN(n639) );
  XOR2_X2 U1042 ( .A(n1367), .B(n639), .Z(n641) );
  XOR2_X2 U1043 ( .A(n1371), .B(n641), .Z(n1378) );
  NAND2_X2 U1044 ( .A1(n1080), .A2(n1077), .ZN(n643) );
  NAND2_X2 U1045 ( .A1(n1097), .A2(n643), .ZN(n649) );
  INV_X4 U1046 ( .A(n649), .ZN(n1341) );
  INV_X4 U1047 ( .A(n1092), .ZN(n645) );
  XOR2_X2 U1048 ( .A(n645), .B(n1091), .Z(n1340) );
  INV_X4 U1049 ( .A(n1340), .ZN(n651) );
  INV_X4 U1050 ( .A(n1094), .ZN(n648) );
  XOR2_X2 U1051 ( .A(n648), .B(n1093), .Z(n1339) );
  NOR2_X2 U1052 ( .A1(n1340), .A2(n649), .ZN(n650) );
  OAI22_X2 U1053 ( .A1(n1341), .A2(n651), .B1(n1339), .B2(n650), .ZN(n1352) );
  OAI22_X2 U1054 ( .A1(n614), .A2(n717), .B1(n590), .B2(n716), .ZN(n715) );
  OAI22_X2 U1055 ( .A1(U1_C_8_), .A2(n715), .B1(n402), .B2(n652), .ZN(n713) );
  OAI22_X2 U1056 ( .A1(n236), .A2(n238), .B1(n824), .B2(n253), .ZN(n867) );
  INV_X4 U1057 ( .A(n658), .ZN(n875) );
  INV_X4 U1058 ( .A(n867), .ZN(n654) );
  NOR2_X2 U1059 ( .A1(n875), .A2(n654), .ZN(n655) );
  OAI22_X2 U1060 ( .A1(n616), .A2(n430), .B1(n595), .B2(n1442), .ZN(n866) );
  OAI22_X2 U1061 ( .A1(n867), .A2(n658), .B1(n655), .B2(n866), .ZN(n667) );
  OAI22_X2 U1062 ( .A1(n236), .A2(n662), .B1(n659), .B2(n254), .ZN(n670) );
  OAI22_X2 U1063 ( .A1(n665), .A2(n430), .B1(n616), .B2(n1442), .ZN(n671) );
  INV_X4 U1064 ( .A(n671), .ZN(n679) );
  INV_X4 U1065 ( .A(n667), .ZN(n711) );
  INV_X4 U1066 ( .A(n713), .ZN(n663) );
  NOR2_X2 U1067 ( .A1(n711), .A2(n663), .ZN(n666) );
  INV_X4 U1068 ( .A(n704), .ZN(n699) );
  OAI22_X2 U1069 ( .A1(n660), .A2(n717), .B1(n614), .B2(n716), .ZN(n690) );
  NAND2_X2 U1070 ( .A1(U1_C_9_), .A2(n690), .ZN(n1004) );
  INV_X4 U1071 ( .A(n670), .ZN(n678) );
  NOR2_X2 U1072 ( .A1(n1548), .A2(n671), .ZN(n677) );
  OAI22_X2 U1073 ( .A1(n661), .A2(n679), .B1(n678), .B2(n677), .ZN(n1002) );
  INV_X4 U1074 ( .A(n1002), .ZN(n1014) );
  XOR2_X2 U1075 ( .A(n444), .B(n436), .Z(n689) );
  INV_X4 U1076 ( .A(n694), .ZN(n748) );
  XOR2_X2 U1077 ( .A(n690), .B(U1_C_9_), .Z(n744) );
  OAI22_X2 U1078 ( .A1(n745), .A2(n694), .B1(n693), .B2(n744), .ZN(n1043) );
  INV_X4 U1079 ( .A(n697), .ZN(n702) );
  NOR2_X2 U1080 ( .A1(n702), .A2(n704), .ZN(n695) );
  OAI22_X2 U1081 ( .A1(n699), .A2(n697), .B1(n703), .B2(n695), .ZN(n1470) );
  INV_X4 U1082 ( .A(n705), .ZN(n712) );
  INV_X4 U1083 ( .A(n743), .ZN(n950) );
  OAI22_X2 U1084 ( .A1(n590), .A2(n717), .B1(n574), .B2(n716), .ZN(n818) );
  NAND2_X2 U1085 ( .A1(n718), .A2(n444), .ZN(n719) );
  INV_X4 U1086 ( .A(n790), .ZN(n734) );
  OAI22_X2 U1087 ( .A1(n595), .A2(n430), .B1(n596), .B2(n1442), .ZN(n730) );
  INV_X4 U1088 ( .A(n730), .ZN(n792) );
  NOR2_X2 U1089 ( .A1(n792), .A2(n790), .ZN(n728) );
  OAI22_X2 U1090 ( .A1(n734), .A2(n730), .B1(n728), .B2(n788), .ZN(n737) );
  NAND2_X2 U1091 ( .A1(n736), .A2(n737), .ZN(n859) );
  NAND2_X2 U1092 ( .A1(n865), .A2(n859), .ZN(n741) );
  NAND3_X2 U1093 ( .A1(U1_C_7_), .A2(n738), .A3(n818), .ZN(n858) );
  NAND2_X2 U1094 ( .A1(n741), .A2(n858), .ZN(n952) );
  INV_X4 U1095 ( .A(n952), .ZN(n742) );
  INV_X4 U1096 ( .A(n773), .ZN(n768) );
  NAND2_X2 U1097 ( .A1(n227), .A2(n1494), .ZN(n780) );
  INV_X4 U1098 ( .A(n781), .ZN(n787) );
  NOR2_X2 U1099 ( .A1(n782), .A2(n781), .ZN(n785) );
  OAI22_X2 U1100 ( .A1(n236), .A2(n824), .B1(n819), .B2(n253), .ZN(n877) );
  INV_X4 U1101 ( .A(n877), .ZN(n901) );
  OAI22_X2 U1102 ( .A1(n828), .A2(U1_C_6_), .B1(n385), .B2(n827), .ZN(n894) );
  INV_X4 U1103 ( .A(n894), .ZN(n880) );
  XOR2_X2 U1104 ( .A(n831), .B(n856), .Z(n1491) );
  INV_X4 U1105 ( .A(n1494), .ZN(n832) );
  INV_X4 U1106 ( .A(n902), .ZN(n1496) );
  INV_X4 U1107 ( .A(n856), .ZN(n851) );
  INV_X4 U1108 ( .A(n904), .ZN(n1497) );
  NAND2_X2 U1109 ( .A1(n859), .A2(n858), .ZN(n863) );
  XNOR2_X2 U1110 ( .A(n865), .B(n863), .ZN(n936) );
  NOR2_X2 U1111 ( .A1(n880), .A2(n877), .ZN(n891) );
  NAND2_X2 U1112 ( .A1(n1496), .A2(n1497), .ZN(n906) );
  NOR2_X2 U1113 ( .A1(n916), .A2(n915), .ZN(n933) );
  OAI22_X2 U1114 ( .A1(n277), .A2(n934), .B1(n933), .B2(n917), .ZN(n1501) );
  INV_X4 U1115 ( .A(n938), .ZN(n951) );
  INV_X4 U1116 ( .A(n968), .ZN(n1469) );
  INV_X4 U1117 ( .A(n969), .ZN(n1466) );
  NOR2_X2 U1118 ( .A1(n1469), .A2(n1466), .ZN(n961) );
  NOR2_X2 U1119 ( .A1(n1471), .A2(n1470), .ZN(n1090) );
  INV_X4 U1120 ( .A(n1138), .ZN(n1134) );
  INV_X4 U1121 ( .A(n987), .ZN(n1015) );
  NOR2_X2 U1122 ( .A1(n1002), .A2(n987), .ZN(n1005) );
  OAI22_X2 U1123 ( .A1(n1015), .A2(n1014), .B1(n1005), .B2(n1004), .ZN(n1133)
         );
  INV_X4 U1124 ( .A(n1133), .ZN(n1139) );
  OAI22_X2 U1125 ( .A1(n1044), .A2(n1043), .B1(n1040), .B2(n1019), .ZN(n1106)
         );
  NAND2_X2 U1126 ( .A1(n1471), .A2(n1470), .ZN(n1073) );
  INV_X4 U1127 ( .A(n1140), .ZN(n1475) );
  XOR2_X2 U1128 ( .A(n1129), .B(n1128), .Z(n1131) );
  XNOR2_X2 U1129 ( .A(n1131), .B(n1130), .ZN(n1155) );
  INV_X4 U1130 ( .A(n1141), .ZN(n1147) );
  NOR2_X2 U1131 ( .A1(n1134), .A2(n1133), .ZN(n1137) );
  INV_X4 U1132 ( .A(n1135), .ZN(n1136) );
  OAI22_X2 U1133 ( .A1(n1139), .A2(n1138), .B1(n1137), .B2(n1136), .ZN(n1146)
         );
  INV_X4 U1134 ( .A(n1146), .ZN(n1142) );
  NOR2_X2 U1135 ( .A1(n1142), .A2(n1141), .ZN(n1145) );
  INV_X4 U1136 ( .A(n1143), .ZN(n1144) );
  OAI22_X2 U1137 ( .A1(n1147), .A2(n1146), .B1(n1145), .B2(n1144), .ZN(n1158)
         );
  INV_X4 U1138 ( .A(n1158), .ZN(n1480) );
  XOR2_X2 U1139 ( .A(n427), .B(in_b_mac[11]), .Z(n1454) );
  XOR2_X2 U1140 ( .A(n1457), .B(n754), .Z(n1149) );
  XNOR2_X2 U1141 ( .A(n1149), .B(n751), .ZN(n1172) );
  INV_X4 U1142 ( .A(n674), .ZN(n1150) );
  XOR2_X2 U1143 ( .A(n1150), .B(n675), .Z(n1162) );
  INV_X4 U1144 ( .A(n1153), .ZN(n1504) );
  XNOR2_X2 U1145 ( .A(n684), .B(n686), .ZN(n1152) );
  XNOR2_X2 U1146 ( .A(n1152), .B(n1151), .ZN(n1154) );
  INV_X4 U1147 ( .A(n1154), .ZN(n1503) );
  NOR2_X2 U1148 ( .A1(n1154), .A2(n1153), .ZN(n1156) );
  INV_X4 U1149 ( .A(n1160), .ZN(n1164) );
  OAI22_X2 U1150 ( .A1(n1164), .A2(n1163), .B1(n1162), .B2(n1161), .ZN(n1176)
         );
  INV_X4 U1151 ( .A(n1176), .ZN(n1483) );
  INV_X4 U1152 ( .A(n1167), .ZN(n1170) );
  NOR2_X2 U1153 ( .A1(n1167), .A2(n1166), .ZN(n1169) );
  OAI22_X2 U1154 ( .A1(n1171), .A2(n1170), .B1(n1169), .B2(n1168), .ZN(n1186)
         );
  OAI22_X2 U1155 ( .A1(n673), .A2(n672), .B1(n750), .B2(n1172), .ZN(n1188) );
  INV_X4 U1156 ( .A(n1188), .ZN(n1185) );
  INV_X4 U1157 ( .A(n1178), .ZN(n1183) );
  NAND2_X2 U1160 ( .A1(n1505), .A2(n707), .ZN(n1174) );
  NAND2_X2 U1164 ( .A1(n706), .A2(n1174), .ZN(n1182) );
  INV_X4 U1167 ( .A(n1182), .ZN(n1177) );
  NOR2_X2 U1168 ( .A1(n1178), .A2(n1177), .ZN(n1181) );
  INV_X4 U1169 ( .A(n1179), .ZN(n1180) );
  OAI22_X2 U1170 ( .A1(n1183), .A2(n1182), .B1(n1181), .B2(n1180), .ZN(n1489)
         );
  INV_X4 U1171 ( .A(n340), .ZN(n1197) );
  INV_X4 U1172 ( .A(n343), .ZN(n1184) );
  NOR2_X2 U1173 ( .A1(n1185), .A2(n1184), .ZN(n1187) );
  OAI22_X2 U1174 ( .A1(n343), .A2(n1188), .B1(n1187), .B2(n1186), .ZN(n1196)
         );
  INV_X4 U1175 ( .A(n1196), .ZN(n1192) );
  INV_X4 U1176 ( .A(n1489), .ZN(n1189) );
  NOR2_X2 U1177 ( .A1(n340), .A2(n1192), .ZN(n1195) );
  INV_X4 U1178 ( .A(n1193), .ZN(n1194) );
  OAI22_X2 U1179 ( .A1(n1197), .A2(n1196), .B1(n1195), .B2(n1194), .ZN(n1205)
         );
  INV_X4 U1180 ( .A(n1205), .ZN(n1393) );
  NAND2_X2 U1181 ( .A1(n770), .A2(n1198), .ZN(n1206) );
  XOR2_X2 U1182 ( .A(n1199), .B(n1546), .Z(n1201) );
  XOR2_X2 U1183 ( .A(n1201), .B(n1200), .Z(n762) );
  XOR2_X2 U1184 ( .A(n762), .B(n765), .Z(n1202) );
  XNOR2_X2 U1185 ( .A(n1202), .B(n764), .ZN(n1209) );
  INV_X4 U1186 ( .A(n1209), .ZN(n1207) );
  INV_X4 U1187 ( .A(n1394), .ZN(n1203) );
  OAI22_X2 U1188 ( .A1(n335), .A2(n1205), .B1(n1204), .B2(n1203), .ZN(n1397)
         );
  INV_X4 U1189 ( .A(n1206), .ZN(n1210) );
  NOR2_X2 U1190 ( .A1(n1207), .A2(n1206), .ZN(n1208) );
  OAI22_X2 U1191 ( .A1(n1210), .A2(n1209), .B1(n1208), .B2(n389), .ZN(n1219)
         );
  INV_X4 U1192 ( .A(n1219), .ZN(n1399) );
  NOR2_X2 U1193 ( .A1(n1397), .A2(n1399), .ZN(n1218) );
  XNOR2_X2 U1194 ( .A(n791), .B(n789), .ZN(n1214) );
  XOR2_X2 U1195 ( .A(n1211), .B(n65), .Z(n1213) );
  XOR2_X2 U1196 ( .A(n1213), .B(n1212), .Z(n1517) );
  XNOR2_X2 U1197 ( .A(n1214), .B(n1517), .ZN(n1227) );
  INV_X4 U1198 ( .A(n1227), .ZN(n1221) );
  OR2_X1 U1199 ( .A1(n794), .A2(n1216), .ZN(n1226) );
  INV_X4 U1200 ( .A(n1226), .ZN(n1222) );
  INV_X4 U1201 ( .A(n1398), .ZN(n1217) );
  OAI22_X2 U1202 ( .A1(n1220), .A2(n1219), .B1(n1218), .B2(n1217), .ZN(n1233)
         );
  NOR2_X2 U1203 ( .A1(n1222), .A2(n1221), .ZN(n1225) );
  INV_X4 U1204 ( .A(n1223), .ZN(n1224) );
  OAI22_X2 U1205 ( .A1(n1227), .A2(n1226), .B1(n1225), .B2(n1224), .ZN(n1401)
         );
  INV_X4 U1206 ( .A(n1401), .ZN(n1228) );
  XOR2_X2 U1207 ( .A(n1229), .B(n836), .Z(n1238) );
  XOR2_X2 U1208 ( .A(n1238), .B(n1237), .Z(n1230) );
  INV_X4 U1209 ( .A(n1234), .ZN(n1239) );
  XNOR2_X2 U1210 ( .A(n1230), .B(n1239), .ZN(n1402) );
  INV_X4 U1211 ( .A(n1402), .ZN(n1231) );
  OAI22_X2 U1212 ( .A1(n312), .A2(n1401), .B1(n1232), .B2(n1231), .ZN(n1248)
         );
  INV_X4 U1213 ( .A(n1238), .ZN(n1235) );
  NOR2_X2 U1214 ( .A1(n1235), .A2(n1234), .ZN(n1236) );
  OAI22_X2 U1215 ( .A1(n1239), .A2(n1238), .B1(n1237), .B2(n1236), .ZN(n1247)
         );
  INV_X4 U1216 ( .A(n1247), .ZN(n1405) );
  XOR2_X2 U1217 ( .A(n1240), .B(n879), .Z(n1241) );
  XNOR2_X2 U1218 ( .A(n1241), .B(n878), .ZN(n1249) );
  XOR2_X2 U1219 ( .A(n926), .B(n927), .Z(n1257) );
  XOR2_X2 U1220 ( .A(n1257), .B(n881), .Z(n1251) );
  XOR2_X2 U1221 ( .A(n1249), .B(n1251), .Z(n1244) );
  INV_X4 U1222 ( .A(n1517), .ZN(n1242) );
  OR2_X1 U1223 ( .A1(n884), .A2(n1243), .ZN(n1253) );
  INV_X4 U1224 ( .A(n1253), .ZN(n1250) );
  XNOR2_X2 U1225 ( .A(n1244), .B(n1250), .ZN(n1406) );
  INV_X4 U1226 ( .A(n1406), .ZN(n1245) );
  OAI22_X2 U1227 ( .A1(n313), .A2(n1247), .B1(n1246), .B2(n1245), .ZN(n1265)
         );
  INV_X4 U1228 ( .A(n1249), .ZN(n1254) );
  NOR2_X2 U1229 ( .A1(n1250), .A2(n1249), .ZN(n1252) );
  OAI22_X2 U1230 ( .A1(n1254), .A2(n1253), .B1(n1252), .B2(n1251), .ZN(n1407)
         );
  INV_X4 U1231 ( .A(n1407), .ZN(n1255) );
  INV_X4 U1232 ( .A(n1265), .ZN(n1409) );
  INV_X4 U1233 ( .A(n888), .ZN(n1256) );
  INV_X4 U1234 ( .A(n1257), .ZN(n1258) );
  OAI22_X2 U1235 ( .A1(n883), .A2(n1502), .B1(n925), .B2(n1258), .ZN(n1270) );
  XOR2_X2 U1236 ( .A(n964), .B(n963), .Z(n1441) );
  XOR2_X2 U1237 ( .A(n1259), .B(n1003), .Z(n1261) );
  XOR2_X2 U1238 ( .A(n1261), .B(n1260), .Z(n918) );
  XOR2_X2 U1239 ( .A(n918), .B(n919), .Z(n1267) );
  INV_X4 U1240 ( .A(n1267), .ZN(n1269) );
  XOR2_X2 U1241 ( .A(n219), .B(n1269), .Z(n1262) );
  XOR2_X2 U1242 ( .A(n1270), .B(n1262), .Z(n1408) );
  INV_X4 U1243 ( .A(n1408), .ZN(n1263) );
  OAI22_X2 U1244 ( .A1(n293), .A2(n1407), .B1(n1264), .B2(n1263), .ZN(n1271)
         );
  INV_X4 U1245 ( .A(n1270), .ZN(n1266) );
  NOR2_X2 U1246 ( .A1(n1267), .A2(n1266), .ZN(n1268) );
  OAI22_X2 U1247 ( .A1(n1270), .A2(n1269), .B1(n219), .B2(n1268), .ZN(n1279)
         );
  INV_X4 U1248 ( .A(n1279), .ZN(n1413) );
  NOR2_X2 U1249 ( .A1(n1271), .A2(n1413), .ZN(n1278) );
  NAND2_X2 U1250 ( .A1(n1515), .A2(n924), .ZN(n1272) );
  NAND2_X2 U1251 ( .A1(n962), .A2(n1272), .ZN(n1283) );
  INV_X4 U1252 ( .A(n958), .ZN(n1273) );
  XOR2_X2 U1253 ( .A(n957), .B(n954), .Z(n1275) );
  INV_X4 U1254 ( .A(n956), .ZN(n1274) );
  XNOR2_X2 U1255 ( .A(n1275), .B(n1274), .ZN(n1280) );
  INV_X4 U1256 ( .A(n1280), .ZN(n1284) );
  XOR2_X2 U1257 ( .A(n222), .B(n1284), .Z(n1276) );
  XOR2_X2 U1258 ( .A(n1283), .B(n1276), .Z(n1412) );
  INV_X4 U1259 ( .A(n1412), .ZN(n1277) );
  INV_X4 U1260 ( .A(n1283), .ZN(n1281) );
  NOR2_X2 U1261 ( .A1(n1281), .A2(n1280), .ZN(n1282) );
  OAI22_X2 U1262 ( .A1(n1284), .A2(n1283), .B1(n1282), .B2(n222), .ZN(n1417)
         );
  INV_X4 U1263 ( .A(n1417), .ZN(n1285) );
  NAND2_X2 U1264 ( .A1(n1518), .A2(n996), .ZN(n1286) );
  NAND2_X2 U1265 ( .A1(n995), .A2(n1286), .ZN(n1295) );
  INV_X4 U1266 ( .A(n991), .ZN(n1287) );
  INV_X4 U1267 ( .A(n988), .ZN(n1288) );
  XOR2_X2 U1268 ( .A(n1288), .B(n989), .Z(n1296) );
  INV_X4 U1269 ( .A(n1296), .ZN(n1292) );
  XOR2_X2 U1270 ( .A(n223), .B(n1292), .Z(n1289) );
  XOR2_X2 U1271 ( .A(n1295), .B(n1289), .Z(n1415) );
  INV_X4 U1272 ( .A(n1295), .ZN(n1293) );
  NOR2_X2 U1273 ( .A1(n1293), .A2(n1292), .ZN(n1294) );
  OAI22_X2 U1274 ( .A1(n1296), .A2(n1295), .B1(n1294), .B2(n223), .ZN(n1421)
         );
  INV_X4 U1275 ( .A(n1421), .ZN(n1297) );
  INV_X4 U1276 ( .A(n1021), .ZN(n1298) );
  XOR2_X2 U1277 ( .A(n1298), .B(n1020), .Z(n1305) );
  INV_X4 U1278 ( .A(n1024), .ZN(n1299) );
  XOR2_X2 U1279 ( .A(n1299), .B(n1025), .Z(n1307) );
  XOR2_X2 U1280 ( .A(n1305), .B(n1307), .Z(n1301) );
  NAND2_X2 U1281 ( .A1(n994), .A2(n993), .ZN(n1300) );
  NAND2_X2 U1282 ( .A1(n1028), .A2(n1300), .ZN(n1304) );
  INV_X4 U1283 ( .A(n1304), .ZN(n1309) );
  XNOR2_X2 U1284 ( .A(n1301), .B(n1309), .ZN(n1419) );
  OAI22_X2 U1285 ( .A1(n1303), .A2(n1421), .B1(n1302), .B2(n1419), .ZN(n1316)
         );
  INV_X4 U1286 ( .A(n1305), .ZN(n1308) );
  NOR2_X2 U1287 ( .A1(n1305), .A2(n1304), .ZN(n1306) );
  OAI22_X2 U1288 ( .A1(n1309), .A2(n1308), .B1(n1307), .B2(n1306), .ZN(n1424)
         );
  NAND2_X2 U1289 ( .A1(n1027), .A2(n1026), .ZN(n1310) );
  NAND2_X2 U1290 ( .A1(n1049), .A2(n1310), .ZN(n1317) );
  INV_X4 U1291 ( .A(n1045), .ZN(n1311) );
  XOR2_X2 U1292 ( .A(n1311), .B(n1046), .Z(n1319) );
  INV_X4 U1293 ( .A(n1319), .ZN(n1322) );
  NAND2_X2 U1294 ( .A1(n1022), .A2(n1021), .ZN(n1312) );
  NAND2_X2 U1295 ( .A1(n1067), .A2(n1312), .ZN(n1318) );
  INV_X4 U1296 ( .A(n1318), .ZN(n1323) );
  XOR2_X2 U1297 ( .A(n1322), .B(n1323), .Z(n1313) );
  XOR2_X2 U1298 ( .A(n1317), .B(n1313), .Z(n1423) );
  INV_X4 U1299 ( .A(n1424), .ZN(n1314) );
  INV_X4 U1300 ( .A(n1317), .ZN(n1321) );
  NOR2_X2 U1301 ( .A1(n1319), .A2(n1318), .ZN(n1320) );
  OAI22_X2 U1302 ( .A1(n1323), .A2(n1322), .B1(n1321), .B2(n1320), .ZN(n1329)
         );
  INV_X4 U1303 ( .A(n1329), .ZN(n1429) );
  INV_X4 U1304 ( .A(n1077), .ZN(n1324) );
  XOR2_X2 U1305 ( .A(n1324), .B(n1078), .Z(n1333) );
  INV_X4 U1306 ( .A(n1074), .ZN(n1325) );
  XOR2_X2 U1307 ( .A(n1325), .B(n1075), .Z(n1332) );
  INV_X4 U1308 ( .A(n1332), .ZN(n1337) );
  XOR2_X2 U1309 ( .A(n1333), .B(n1337), .Z(n1327) );
  NOR2_X2 U1310 ( .A1(n1048), .A2(n1047), .ZN(n1326) );
  OR2_X1 U1311 ( .A1(n1081), .A2(n1326), .ZN(n1336) );
  INV_X4 U1312 ( .A(n1336), .ZN(n1331) );
  XOR2_X2 U1313 ( .A(n1327), .B(n1331), .Z(n1427) );
  OAI22_X2 U1314 ( .A1(n1330), .A2(n1329), .B1(n1328), .B2(n1427), .ZN(n1344)
         );
  NOR2_X2 U1315 ( .A1(n1332), .A2(n1331), .ZN(n1335) );
  INV_X4 U1316 ( .A(n1333), .ZN(n1334) );
  OAI22_X2 U1317 ( .A1(n1337), .A2(n1336), .B1(n1335), .B2(n1334), .ZN(n1432)
         );
  INV_X4 U1318 ( .A(n1432), .ZN(n1338) );
  XOR2_X2 U1319 ( .A(n1340), .B(n1339), .Z(n1342) );
  XNOR2_X2 U1320 ( .A(n1342), .B(n1341), .ZN(n1431) );
  INV_X4 U1321 ( .A(n1352), .ZN(n1434) );
  INV_X4 U1322 ( .A(n1107), .ZN(n1345) );
  XOR2_X2 U1323 ( .A(n1345), .B(n1108), .Z(n1353) );
  INV_X4 U1324 ( .A(n1096), .ZN(n1532) );
  NOR2_X2 U1325 ( .A1(n1094), .A2(n1532), .ZN(n1346) );
  OR2_X1 U1326 ( .A1(n1110), .A2(n1346), .ZN(n1355) );
  XOR2_X2 U1327 ( .A(n1353), .B(n1355), .Z(n1348) );
  NAND2_X2 U1328 ( .A1(n1092), .A2(U1_C_25_), .ZN(n1347) );
  NAND2_X2 U1329 ( .A1(n1116), .A2(n1347), .ZN(n1357) );
  INV_X4 U1330 ( .A(n1357), .ZN(n1354) );
  XNOR2_X2 U1331 ( .A(n1348), .B(n1354), .ZN(n1435) );
  INV_X4 U1332 ( .A(n1435), .ZN(n1349) );
  OAI22_X2 U1333 ( .A1(n1352), .A2(n292), .B1(n1350), .B2(n1349), .ZN(n1365)
         );
  INV_X4 U1334 ( .A(n1353), .ZN(n1358) );
  NOR2_X2 U1335 ( .A1(n1354), .A2(n1353), .ZN(n1356) );
  INV_X4 U1336 ( .A(n1438), .ZN(n1359) );
  INV_X4 U1337 ( .A(n1365), .ZN(n1440) );
  NOR2_X2 U1338 ( .A1(n1440), .A2(n1359), .ZN(n1364) );
  XOR2_X2 U1339 ( .A(n1360), .B(n224), .Z(n1362) );
  XOR2_X2 U1340 ( .A(n1362), .B(n1361), .Z(n1439) );
  NOR2_X2 U1341 ( .A1(n208), .A2(n215), .ZN(U6_Z_29) );
  INV_X4 U1342 ( .A(n1371), .ZN(n1368) );
  NOR2_X2 U1343 ( .A1(n1368), .A2(n1367), .ZN(n1370) );
  OAI22_X2 U1344 ( .A1(n4), .A2(n1371), .B1(n1370), .B2(n1369), .ZN(n1384) );
  NAND2_X2 U1345 ( .A1(n360), .A2(n361), .ZN(n1373) );
  INV_X4 U1346 ( .A(n362), .ZN(n1372) );
  NAND2_X2 U1347 ( .A1(n1373), .A2(n1372), .ZN(n1389) );
  XOR2_X2 U1348 ( .A(U1_C_30_), .B(n1367), .Z(n1374) );
  XOR2_X2 U1349 ( .A(n1389), .B(n1374), .Z(n1382) );
  INV_X4 U1350 ( .A(n1382), .ZN(n1387) );
  INV_X4 U1351 ( .A(n1379), .ZN(n1376) );
  INV_X4 U1352 ( .A(n1386), .ZN(n1383) );
  NOR2_X2 U1353 ( .A1(n208), .A2(n396), .ZN(U6_Z_30) );
  OAI22_X2 U1354 ( .A1(n1387), .A2(n308), .B1(n1385), .B2(n1384), .ZN(n1392)
         );
  NOR2_X2 U1355 ( .A1(n4), .A2(n1388), .ZN(n1390) );
  OAI22_X2 U1356 ( .A1(U1_C_30_), .A2(n1367), .B1(n1390), .B2(n1389), .ZN(
        n1391) );
  XOR2_X2 U1357 ( .A(n1394), .B(n1393), .Z(n1396) );
  XNOR2_X2 U1358 ( .A(n1400), .B(n1399), .ZN(n257) );
  XNOR2_X2 U1359 ( .A(n1402), .B(n1401), .ZN(n1404) );
  XNOR2_X2 U1360 ( .A(n1408), .B(n1407), .ZN(n1410) );
  XOR2_X2 U1361 ( .A(n1412), .B(n1411), .Z(n1414) );
  XOR2_X2 U1362 ( .A(n1414), .B(n1413), .Z(n249) );
  XNOR2_X2 U1363 ( .A(n1418), .B(n1417), .ZN(n248) );
  XNOR2_X2 U1364 ( .A(n1422), .B(n1421), .ZN(n247) );
  XNOR2_X2 U1365 ( .A(n1430), .B(n1429), .ZN(n245) );
  XOR2_X2 U1366 ( .A(n1432), .B(n1431), .Z(n1433) );
  XOR2_X2 U1367 ( .A(n1435), .B(n1434), .Z(n1437) );
  INV_X4 U1368 ( .A(n1441), .ZN(n922) );
  INV_X4 U1369 ( .A(n1518), .ZN(n960) );
  INV_X4 U1370 ( .A(n996), .ZN(n1520) );
  XOR2_X2 U1371 ( .A(n939), .B(n1443), .Z(n937) );
  INV_X4 U1372 ( .A(n848), .ZN(n1527) );
  OAI22_X2 U1373 ( .A1(n1448), .A2(n1453), .B1(n862), .B2(n864), .ZN(n847) );
  XOR2_X2 U1374 ( .A(n352), .B(in_b_mac[12]), .Z(n1455) );
  INV_X4 U1375 ( .A(n1461), .ZN(n1452) );
  NOR2_X2 U1376 ( .A1(n1452), .A2(n1451), .ZN(n1531) );
  INV_X4 U1377 ( .A(n1508), .ZN(n845) );
  OAI22_X2 U1378 ( .A1(n1456), .A2(n1462), .B1(n777), .B2(n779), .ZN(n774) );
  INV_X4 U1379 ( .A(n1457), .ZN(n1459) );
  NOR2_X2 U1380 ( .A1(n1459), .A2(n1458), .ZN(n1538) );
  NAND2_X2 U1381 ( .A1(U1_C_13_), .A2(n1460), .ZN(n739) );
  INV_X4 U1382 ( .A(n739), .ZN(n1507) );
  INV_X4 U1383 ( .A(n808), .ZN(n1537) );
  XOR2_X2 U1384 ( .A(n1461), .B(n806), .Z(n804) );
  INV_X4 U1385 ( .A(n1463), .ZN(n1465) );
  NOR2_X2 U1386 ( .A1(n1465), .A2(n1464), .ZN(n1543) );
  XOR2_X2 U1387 ( .A(n1469), .B(n1468), .Z(n283) );
  XNOR2_X2 U1388 ( .A(n1476), .B(n1475), .ZN(n1478) );
  XOR2_X2 U1389 ( .A(n1480), .B(n1479), .Z(n1481) );
  XNOR2_X2 U1390 ( .A(n1484), .B(n1483), .ZN(n1486) );
  INV_X4 U1391 ( .A(n1487), .ZN(n1488) );
  INV_X4 U1392 ( .A(n799), .ZN(n1506) );
  INV_X4 U1393 ( .A(n895), .ZN(n1510) );
  INV_X4 U1394 ( .A(n789), .ZN(n1511) );
  INV_X4 U1395 ( .A(n885), .ZN(n1512) );
  INV_X4 U1396 ( .A(n897), .ZN(n1514) );
  INV_X4 U1397 ( .A(n930), .ZN(n1516) );
  INV_X4 U1398 ( .A(n1038), .ZN(n1519) );
  INV_X4 U1399 ( .A(n1053), .ZN(n1521) );
  INV_X4 U1400 ( .A(n1054), .ZN(n1522) );
  INV_X4 U1401 ( .A(n1087), .ZN(n1523) );
  INV_X4 U1402 ( .A(n1112), .ZN(n1524) );
  INV_X4 U1403 ( .A(n1085), .ZN(n1525) );
  INV_X4 U1404 ( .A(n1083), .ZN(n1528) );
  INV_X4 U1405 ( .A(n1061), .ZN(n1529) );
  INV_X4 U1406 ( .A(n843), .ZN(n1530) );
  INV_X4 U1407 ( .A(n1070), .ZN(n1533) );
  INV_X4 U1408 ( .A(n1057), .ZN(n1534) );
  INV_X4 U1409 ( .A(n1008), .ZN(n1535) );
  INV_X4 U1410 ( .A(n941), .ZN(n1536) );
  INV_X4 U1411 ( .A(n1101), .ZN(n1539) );
  INV_X4 U1412 ( .A(n1031), .ZN(n1540) );
  INV_X4 U1413 ( .A(n932), .ZN(n1541) );
  INV_X4 U1414 ( .A(n947), .ZN(n1542) );
  INV_X4 U1415 ( .A(n982), .ZN(n1544) );
  INV_X4 U1416 ( .A(n870), .ZN(n1545) );
  INV_X4 U1417 ( .A(n903), .ZN(n1546) );
  INV_X4 U1418 ( .A(n811), .ZN(n1547) );
  INV_X4 U1419 ( .A(n709), .ZN(n1549) );
  INV_X4 U1420 ( .A(n642), .ZN(n1550) );
endmodule


module macopertion_m ( in_z_mac, in_m_mac, sendz_count, clk, minm );
  input [15:0] in_z_mac;
  input [15:0] in_m_mac;
  input [5:0] sendz_count;
  output [15:0] minm;
  input clk;
  wire   U6_Z_0, U6_Z_1, U6_Z_2, U6_Z_3, U6_Z_4, U6_Z_5, U6_Z_6, U6_Z_7,
         U6_Z_8, U6_Z_9, U6_Z_10, U6_Z_11, U6_Z_12, U6_Z_13, U6_Z_14, U6_Z_15,
         U6_Z_16, U6_Z_17, U6_Z_18, U6_Z_19, U6_Z_20, U6_Z_21, U6_Z_22,
         U6_Z_23, U6_Z_24, U6_Z_25, U6_Z_26, U6_Z_27, U6_Z_28, U6_Z_29,
         U6_Z_30, U5_Z_0, U5_Z_1, U5_Z_2, U5_Z_3, U5_Z_4, U5_Z_5, U5_Z_6,
         U5_Z_7, U5_Z_8, U5_Z_9, U5_Z_10, U5_Z_11, U5_Z_12, U5_Z_13, U5_Z_14,
         U1_C_31_, U1_C_30_, U1_C_28_, U1_C_26_, U1_C_24_, U1_C_22_, U1_C_20_,
         U1_C_18_, U1_C_16_, U1_C_15_, U1_C_14_, U1_C_13_, U1_C_12_, U1_C_11_,
         U1_C_10_, U1_C_9_, U1_C_8_, U1_C_7_, U1_C_6_, U1_C_5_, U1_C_4_,
         U1_C_3_, U1_C_2_, U1_C_1_, U1_C_0_, U1_C_17_, U1_C_21_, U1_C_23_,
         U1_C_25_, U1_C_27_, n4, n12, n18, n29, n41, n52, n65, n208, n209,
         n212, n217, n242, n243, n244, n245, n247, n248, n249, n250, n255,
         n256, n257, n258, n259, n264, n269, n274, n279, n283, n294, n361,
         n363, n367, n368, n369, n560, n575, n591, n596, n597, n614, n615,
         n617, n622, n624, n625, n636, n641, n643, n645, n647, n648, n654,
         n657, n658, n661, n662, n665, n666, n673, n674, n675, n676, n677,
         n685, n687, n689, n692, n693, n697, n699, n701, n702, n707, n708,
         n709, n710, n711, n715, n721, n722, n723, n725, n726, n727, n730,
         n731, n732, n733, n734, n736, n740, n741, n747, n748, n751, n752,
         n755, n757, n758, n761, n763, n765, n766, n767, n770, n771, n774,
         n775, n776, n777, n778, n779, n780, n784, n790, n792, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n806, n807,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n821,
         n822, n823, n824, n826, n827, n830, n831, n834, n836, n837, n838,
         n839, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n853, n855, n861, n862, n863, n865, n869, n870, n871, n872, n873,
         n874, n875, n877, n879, n880, n882, n884, n885, n886, n887, n888,
         n889, n890, n891, n893, n894, n896, n897, n898, n899, n900, n901,
         n904, n906, n908, n909, n910, n911, n912, n913, n914, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n936, n938, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n955, n957, n958, n959, n960, n961, n963,
         n964, n965, n966, n967, n968, n971, n972, n973, n974, n976, n977,
         n979, n980, n981, n983, n984, n985, n987, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1004,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1017, n1019,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1042, n1043, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
         n1117, n1118, n1120, n1121, n1122, n1123, n1124, n1125, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n210, n211, n213, n214, n215, n216, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n246, n251,
         n252, n253, n254, n260, n261, n262, n263, n265, n266, n267, n268,
         n270, n271, n272, n273, n275, n276, n277, n278, n280, n281, n282,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n362,
         n364, n365, n366, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n592, n593, n594, n595, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n616, n618, n619, n620, n621, n623, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n637, n638, n639, n640, n642, n644,
         n646, n649, n650, n651, n652, n653, n655, n656, n659, n660, n663,
         n664, n667, n668, n669, n670, n671, n672, n678, n679, n680, n681,
         n682, n683, n684, n686, n688, n690, n691, n694, n695, n696, n698,
         n700, n703, n704, n705, n706, n712, n713, n714, n716, n717, n718,
         n719, n720, n724, n728, n729, n735, n737, n738, n739, n742, n743,
         n744, n745, n746, n749, n750, n753, n754, n756, n759, n760, n762,
         n764, n768, n769, n772, n773, n781, n782, n783, n785, n786, n787,
         n788, n789, n791, n793, n805, n808, n819, n820, n825, n828, n829,
         n832, n833, n835, n840, n851, n852, n854, n856, n857, n858, n859,
         n860, n864, n866, n867, n868, n876, n878, n881, n883, n892, n895,
         n902, n903, n905, n907, n915, n916, n917, n918, n934, n935, n937,
         n939, n951, n952, n953, n954, n956, n962, n969, n970, n975, n978,
         n982, n986, n988, n1003, n1005, n1006, n1015, n1016, n1018, n1020,
         n1041, n1044, n1045, n1074, n1091, n1107, n1119, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
         n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
         n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
         n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
         n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
         n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
         n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
         n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
         n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
         n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
         n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
         n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
         n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
         n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
         n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
         n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
         n1569, n1570, n1571, n1572, n1573, n1574, n1575;
  assign minm[15] = 1'b0;

  NOR2_X2 U6 ( .A1(n208), .A2(n209), .ZN(U6_Z_9) );
  NOR2_X2 U9 ( .A1(n208), .A2(n212), .ZN(U6_Z_8) );
  NOR2_X2 U12 ( .A1(n208), .A2(n217), .ZN(U6_Z_7) );
  NOR2_X2 U29 ( .A1(n208), .A2(n242), .ZN(U6_Z_28) );
  NOR2_X2 U30 ( .A1(n208), .A2(n243), .ZN(U6_Z_27) );
  NOR2_X2 U31 ( .A1(n208), .A2(n244), .ZN(U6_Z_26) );
  NOR2_X2 U32 ( .A1(n208), .A2(n245), .ZN(U6_Z_25) );
  NOR2_X2 U33 ( .A1(n208), .A2(n223), .ZN(U6_Z_24) );
  NOR2_X2 U34 ( .A1(n208), .A2(n247), .ZN(U6_Z_23) );
  NOR2_X2 U35 ( .A1(n208), .A2(n248), .ZN(U6_Z_22) );
  NOR2_X2 U36 ( .A1(n208), .A2(n249), .ZN(U6_Z_21) );
  NOR2_X2 U37 ( .A1(n208), .A2(n250), .ZN(U6_Z_20) );
  NOR2_X2 U41 ( .A1(n208), .A2(n255), .ZN(U6_Z_19) );
  NOR2_X2 U42 ( .A1(n208), .A2(n256), .ZN(U6_Z_18) );
  NOR2_X2 U43 ( .A1(n208), .A2(n257), .ZN(U6_Z_17) );
  NOR2_X2 U44 ( .A1(n208), .A2(n258), .ZN(U6_Z_16) );
  NOR2_X2 U45 ( .A1(n208), .A2(n259), .ZN(U6_Z_15) );
  NOR2_X2 U48 ( .A1(n208), .A2(n264), .ZN(U6_Z_14) );
  NOR2_X2 U51 ( .A1(n208), .A2(n269), .ZN(U6_Z_13) );
  NOR2_X2 U54 ( .A1(n208), .A2(n274), .ZN(U6_Z_12) );
  NOR2_X2 U57 ( .A1(n208), .A2(n279), .ZN(U6_Z_11) );
  NOR2_X2 U60 ( .A1(n208), .A2(n283), .ZN(U6_Z_10) );
  XOR2_X2 U132 ( .A(in_m_mac[15]), .B(n1575), .Z(n363) );
  XOR2_X2 U336 ( .A(n1572), .B(n459), .Z(n597) );
  OAI22_X2 U421 ( .A1(n468), .A2(n692), .B1(n641), .B2(n643), .ZN(n636) );
  XNOR2_X2 U440 ( .A(n709), .B(n1568), .ZN(n675) );
  XOR2_X2 U441 ( .A(n710), .B(n711), .Z(n709) );
  OAI22_X2 U457 ( .A1(n466), .A2(n725), .B1(n726), .B2(n722), .ZN(n654) );
  XNOR2_X2 U466 ( .A(n732), .B(n733), .ZN(n731) );
  OAI22_X2 U486 ( .A1(n466), .A2(n757), .B1(n725), .B2(n722), .ZN(n687) );
  XOR2_X2 U495 ( .A(in_m_mac[5]), .B(n1572), .Z(n727) );
  XOR2_X2 U513 ( .A(n775), .B(n776), .Z(n774) );
  XNOR2_X2 U516 ( .A(n778), .B(n779), .ZN(n702) );
  XOR2_X2 U530 ( .A(n796), .B(n797), .Z(n767) );
  XOR2_X2 U531 ( .A(n798), .B(n799), .Z(n797) );
  XOR2_X2 U534 ( .A(n801), .B(n802), .Z(n730) );
  XOR2_X2 U535 ( .A(n803), .B(n804), .Z(n802) );
  OAI22_X2 U542 ( .A1(n464), .A2(n813), .B1(n814), .B2(n815), .ZN(n711) );
  XOR2_X2 U555 ( .A(in_m_mac[6]), .B(n1572), .Z(n761) );
  OAI22_X2 U556 ( .A1(n466), .A2(n822), .B1(n757), .B2(n722), .ZN(n755) );
  OAI22_X2 U562 ( .A1(n464), .A2(n826), .B1(n813), .B2(n815), .ZN(n780) );
  OAI22_X2 U564 ( .A1(n466), .A2(n827), .B1(n822), .B2(n722), .ZN(n778) );
  XOR2_X2 U584 ( .A(n838), .B(n839), .Z(n837) );
  XNOR2_X2 U589 ( .A(n1530), .B(n847), .ZN(n794) );
  XNOR2_X2 U590 ( .A(n848), .B(n849), .ZN(n847) );
  XNOR2_X2 U595 ( .A(n1535), .B(n853), .ZN(n766) );
  XNOR2_X2 U596 ( .A(n446), .B(n855), .ZN(n853) );
  OAI22_X2 U604 ( .A1(n798), .A2(n799), .B1(n862), .B2(n796), .ZN(n844) );
  OAI22_X2 U612 ( .A1(n466), .A2(n870), .B1(n827), .B2(n722), .ZN(n806) );
  OAI22_X2 U616 ( .A1(n465), .A2(n872), .B1(n873), .B2(n361), .ZN(n803) );
  OAI22_X2 U620 ( .A1(n464), .A2(n875), .B1(n826), .B2(n815), .ZN(n804) );
  XOR2_X2 U621 ( .A(n320), .B(n1574), .Z(n826) );
  XOR2_X2 U627 ( .A(n1523), .B(n884), .Z(n882) );
  XNOR2_X2 U630 ( .A(n886), .B(n887), .ZN(n841) );
  XOR2_X2 U631 ( .A(n888), .B(n889), .Z(n887) );
  OAI22_X2 U636 ( .A1(n465), .A2(n893), .B1(n872), .B2(n361), .ZN(n865) );
  OAI22_X2 U638 ( .A1(n464), .A2(n894), .B1(n875), .B2(n815), .ZN(n863) );
  OAI22_X2 U653 ( .A1(n466), .A2(n906), .B1(n870), .B2(n722), .ZN(n904) );
  XOR2_X2 U654 ( .A(in_m_mac[5]), .B(n1573), .Z(n870) );
  XNOR2_X2 U660 ( .A(n909), .B(n910), .ZN(n792) );
  XOR2_X2 U661 ( .A(n911), .B(n912), .Z(n910) );
  XOR2_X2 U662 ( .A(n1534), .B(n913), .Z(n790) );
  XNOR2_X2 U663 ( .A(n914), .B(n1563), .ZN(n913) );
  XOR2_X2 U669 ( .A(n921), .B(n922), .Z(n920) );
  XOR2_X2 U671 ( .A(n1536), .B(n925), .Z(n924) );
  XOR2_X2 U674 ( .A(n929), .B(n930), .Z(n928) );
  XNOR2_X2 U677 ( .A(n932), .B(n933), .ZN(n839) );
  XOR2_X2 U678 ( .A(U1_C_18_), .B(n65), .Z(n932) );
  XOR2_X2 U681 ( .A(n938), .B(n1565), .Z(n838) );
  OAI22_X2 U687 ( .A1(n465), .A2(n943), .B1(n893), .B2(n361), .ZN(n911) );
  XOR2_X2 U688 ( .A(n320), .B(n1575), .Z(n893) );
  OAI22_X2 U689 ( .A1(n464), .A2(n944), .B1(n894), .B2(n815), .ZN(n909) );
  OAI22_X2 U694 ( .A1(n466), .A2(n949), .B1(n906), .B2(n722), .ZN(n914) );
  XOR2_X2 U695 ( .A(in_m_mac[6]), .B(n1573), .Z(n906) );
  NOR2_X2 U696 ( .A1(n899), .A2(U1_C_16_), .ZN(n900) );
  XOR2_X2 U698 ( .A(in_m_mac[9]), .B(n1572), .Z(n861) );
  XOR2_X2 U699 ( .A(in_m_mac[10]), .B(n1572), .Z(n946) );
  XOR2_X2 U713 ( .A(n961), .B(n1541), .Z(n960) );
  XNOR2_X2 U717 ( .A(n966), .B(n967), .ZN(n964) );
  XNOR2_X2 U722 ( .A(n971), .B(n972), .ZN(n880) );
  XOR2_X2 U723 ( .A(n973), .B(n974), .Z(n972) );
  OAI22_X2 U726 ( .A1(n464), .A2(n976), .B1(n944), .B2(n815), .ZN(n936) );
  XOR2_X2 U727 ( .A(in_m_mac[5]), .B(n1574), .Z(n944) );
  XOR2_X2 U729 ( .A(in_m_mac[11]), .B(n1572), .Z(n945) );
  OAI22_X2 U740 ( .A1(n465), .A2(n984), .B1(n943), .B2(n361), .ZN(n940) );
  OAI22_X2 U749 ( .A1(n464), .A2(n987), .B1(n976), .B2(n815), .ZN(n930) );
  XOR2_X2 U750 ( .A(in_m_mac[6]), .B(n1574), .Z(n976) );
  XOR2_X2 U754 ( .A(n991), .B(n1550), .Z(n990) );
  XOR2_X2 U756 ( .A(n994), .B(n995), .Z(n993) );
  XOR2_X2 U759 ( .A(n998), .B(n999), .Z(n959) );
  XOR2_X2 U760 ( .A(n1000), .B(n1001), .Z(n999) );
  OAI22_X2 U761 ( .A1(n921), .A2(n922), .B1(n1002), .B2(n919), .ZN(n997) );
  XOR2_X2 U764 ( .A(n1007), .B(n1008), .Z(n922) );
  XNOR2_X2 U765 ( .A(U1_C_20_), .B(n609), .ZN(n1007) );
  OAI22_X2 U768 ( .A1(n465), .A2(n1010), .B1(n984), .B2(n361), .ZN(n973) );
  OAI22_X2 U770 ( .A1(n466), .A2(n1011), .B1(n985), .B2(n722), .ZN(n971) );
  OAI22_X2 U776 ( .A1(n465), .A2(n1014), .B1(n1010), .B2(n361), .ZN(n967) );
  XOR2_X2 U777 ( .A(in_m_mac[5]), .B(n1575), .Z(n1010) );
  XOR2_X2 U781 ( .A(in_m_mac[12]), .B(n1572), .Z(n977) );
  OAI22_X2 U784 ( .A1(n464), .A2(n1019), .B1(n987), .B2(n815), .ZN(n966) );
  XOR2_X2 U785 ( .A(in_m_mac[7]), .B(n1574), .Z(n987) );
  XNOR2_X2 U789 ( .A(n1023), .B(n1024), .ZN(n1021) );
  XOR2_X2 U791 ( .A(n1027), .B(n1028), .Z(n1026) );
  XOR2_X2 U794 ( .A(n1030), .B(n1554), .Z(n992) );
  XOR2_X2 U795 ( .A(U1_C_22_), .B(n41), .Z(n1030) );
  XNOR2_X2 U796 ( .A(n1031), .B(n1032), .ZN(n995) );
  XOR2_X2 U797 ( .A(n1033), .B(n1034), .Z(n1031) );
  XNOR2_X2 U800 ( .A(n1036), .B(n1037), .ZN(n955) );
  XOR2_X2 U801 ( .A(n41), .B(n1038), .Z(n1037) );
  XOR2_X2 U809 ( .A(in_m_mac[13]), .B(n1572), .Z(n1017) );
  OAI22_X2 U810 ( .A1(n466), .A2(n1043), .B1(n1011), .B2(n722), .ZN(n1004) );
  XOR2_X2 U811 ( .A(in_m_mac[9]), .B(n1573), .Z(n1011) );
  XOR2_X2 U819 ( .A(n1048), .B(n1049), .Z(n1047) );
  XOR2_X2 U822 ( .A(n1051), .B(n1052), .Z(n1025) );
  XOR2_X2 U823 ( .A(n29), .B(n1053), .Z(n1052) );
  XOR2_X2 U831 ( .A(in_m_mac[14]), .B(n1572), .Z(n1042) );
  OAI22_X2 U834 ( .A1(n464), .A2(n1059), .B1(n1019), .B2(n815), .ZN(n1000) );
  OAI22_X2 U836 ( .A1(n466), .A2(n1060), .B1(n1043), .B2(n722), .ZN(n998) );
  XOR2_X2 U837 ( .A(in_m_mac[10]), .B(n1573), .Z(n1043) );
  OAI22_X2 U838 ( .A1(n465), .A2(n1061), .B1(n1014), .B2(n361), .ZN(n1001) );
  XOR2_X2 U839 ( .A(in_m_mac[6]), .B(n1575), .Z(n1014) );
  OAI22_X2 U844 ( .A1(n465), .A2(n1065), .B1(n1061), .B2(n361), .ZN(n1034) );
  XOR2_X2 U845 ( .A(in_m_mac[7]), .B(n1575), .Z(n1061) );
  OAI22_X2 U846 ( .A1(n464), .A2(n1066), .B1(n1059), .B2(n815), .ZN(n1032) );
  XOR2_X2 U847 ( .A(in_m_mac[9]), .B(n1574), .Z(n1059) );
  XOR2_X2 U849 ( .A(in_m_mac[15]), .B(n1572), .Z(n1057) );
  OAI22_X2 U855 ( .A1(n465), .A2(n1069), .B1(n1065), .B2(n361), .ZN(n1024) );
  OAI22_X2 U859 ( .A1(n466), .A2(n1072), .B1(n1060), .B2(n722), .ZN(n1071) );
  XOR2_X2 U860 ( .A(in_m_mac[11]), .B(n1573), .Z(n1060) );
  OAI22_X2 U861 ( .A1(n464), .A2(n1073), .B1(n1066), .B2(n815), .ZN(n1023) );
  XOR2_X2 U862 ( .A(in_m_mac[10]), .B(n1574), .Z(n1066) );
  XOR2_X2 U866 ( .A(n18), .B(n1077), .Z(n1076) );
  XOR2_X2 U868 ( .A(n1080), .B(n1081), .Z(n1079) );
  XOR2_X2 U871 ( .A(n1083), .B(n1084), .Z(n1046) );
  XOR2_X2 U872 ( .A(U1_C_24_), .B(n29), .Z(n1083) );
  XNOR2_X2 U873 ( .A(n1085), .B(n1560), .ZN(n1049) );
  XOR2_X2 U874 ( .A(n1086), .B(n1087), .Z(n1085) );
  OAI22_X2 U877 ( .A1(n466), .A2(n1089), .B1(n1072), .B2(n722), .ZN(n1051) );
  XOR2_X2 U878 ( .A(in_m_mac[12]), .B(n1573), .Z(n1072) );
  XOR2_X2 U884 ( .A(U1_C_26_), .B(n18), .Z(n1092) );
  XOR2_X2 U886 ( .A(n1096), .B(n1097), .Z(n1094) );
  OAI22_X2 U891 ( .A1(n466), .A2(n1100), .B1(n1089), .B2(n722), .ZN(n1084) );
  XOR2_X2 U892 ( .A(in_m_mac[13]), .B(n1573), .Z(n1089) );
  OAI22_X2 U895 ( .A1(n464), .A2(n1103), .B1(n1073), .B2(n815), .ZN(n1087) );
  XOR2_X2 U896 ( .A(in_m_mac[11]), .B(n1574), .Z(n1073) );
  OAI22_X2 U897 ( .A1(n465), .A2(n1104), .B1(n1069), .B2(n361), .ZN(n1102) );
  XOR2_X2 U898 ( .A(in_m_mac[9]), .B(n1575), .Z(n1069) );
  OAI22_X2 U904 ( .A1(n465), .A2(n1106), .B1(n1104), .B2(n361), .ZN(n1081) );
  XOR2_X2 U905 ( .A(in_m_mac[10]), .B(n1575), .Z(n1104) );
  XOR2_X2 U909 ( .A(n12), .B(n1110), .Z(n1109) );
  OAI22_X2 U915 ( .A1(n464), .A2(n1114), .B1(n1103), .B2(n815), .ZN(n1075) );
  XOR2_X2 U916 ( .A(in_m_mac[12]), .B(n1574), .Z(n1103) );
  OAI22_X2 U917 ( .A1(n466), .A2(n1112), .B1(n1100), .B2(n722), .ZN(n1077) );
  XOR2_X2 U919 ( .A(in_z_mac[11]), .B(in_z_mac[10]), .Z(n1115) );
  XOR2_X2 U920 ( .A(in_m_mac[14]), .B(n1573), .Z(n1100) );
  XOR2_X2 U921 ( .A(in_m_mac[15]), .B(n1573), .Z(n1112) );
  OAI22_X2 U923 ( .A1(n465), .A2(n1116), .B1(n1106), .B2(n361), .ZN(n1097) );
  XOR2_X2 U924 ( .A(in_m_mac[11]), .B(n1575), .Z(n1106) );
  OAI22_X2 U927 ( .A1(n464), .A2(n1118), .B1(n1114), .B2(n815), .ZN(n1093) );
  XOR2_X2 U928 ( .A(in_m_mac[13]), .B(n1574), .Z(n1114) );
  OAI22_X2 U932 ( .A1(n465), .A2(n369), .B1(n1121), .B2(n361), .ZN(n368) );
  XOR2_X2 U933 ( .A(in_m_mac[14]), .B(n1575), .Z(n369) );
  XOR2_X2 U934 ( .A(U1_C_28_), .B(n12), .Z(n1120) );
  OAI22_X2 U937 ( .A1(n465), .A2(n1121), .B1(n1116), .B2(n361), .ZN(n1108) );
  XOR2_X2 U939 ( .A(in_z_mac[15]), .B(in_z_mac[14]), .Z(n1123) );
  XOR2_X2 U940 ( .A(in_m_mac[12]), .B(n1575), .Z(n1116) );
  XOR2_X2 U941 ( .A(in_m_mac[13]), .B(n1575), .Z(n1121) );
  OAI22_X2 U943 ( .A1(n464), .A2(n1124), .B1(n1118), .B2(n815), .ZN(n1110) );
  XOR2_X2 U944 ( .A(in_m_mac[14]), .B(n1574), .Z(n1118) );
  XOR2_X2 U946 ( .A(in_m_mac[15]), .B(n1574), .Z(n1124) );
  XOR2_X2 U948 ( .A(in_z_mac[13]), .B(in_z_mac[12]), .Z(n1125) );
  OR3_X1 U1149 ( .A1(sendz_count[5]), .A2(sendz_count[4]), .A3(sendz_count[3]), 
        .ZN(n294) );
  OR2_X1 U1159 ( .A1(n459), .A2(n466), .ZN(n721) );
  AND2_X1 U1160 ( .A1(n674), .A2(n673), .ZN(n751) );
  OR2_X1 U1162 ( .A1(n459), .A2(n464), .ZN(n816) );
  AND2_X1 U1163 ( .A1(n799), .A2(n798), .ZN(n862) );
  OR2_X1 U1164 ( .A1(n459), .A2(n465), .ZN(n869) );
  AND2_X1 U1166 ( .A1(n884), .A2(n1523), .ZN(n926) );
  AND2_X1 U1167 ( .A1(n922), .A2(n921), .ZN(n1002) );
  DFF_X2 in_cm_mac_reg_30_ ( .D(U6_Z_30), .CK(clk), .Q(U1_C_30_), .QN(n1405)
         );
  DFF_X2 minm_reg_13_ ( .D(U5_Z_13), .CK(clk), .Q(minm[13]) );
  DFF_X2 minm_reg_12_ ( .D(U5_Z_12), .CK(clk), .Q(minm[12]) );
  DFF_X2 minm_reg_8_ ( .D(U5_Z_8), .CK(clk), .Q(minm[8]) );
  DFF_X2 minm_reg_10_ ( .D(U5_Z_10), .CK(clk), .Q(minm[10]) );
  DFF_X2 minm_reg_9_ ( .D(U5_Z_9), .CK(clk), .Q(minm[9]) );
  DFF_X2 minm_reg_4_ ( .D(U5_Z_4), .CK(clk), .Q(minm[4]) );
  DFF_X2 minm_reg_3_ ( .D(U5_Z_3), .CK(clk), .Q(minm[3]) );
  DFF_X2 minm_reg_14_ ( .D(U5_Z_14), .CK(clk), .Q(minm[14]) );
  DFF_X2 in_cm_mac_reg_26_ ( .D(U6_Z_26), .CK(clk), .Q(U1_C_26_) );
  DFF_X2 in_cm_mac_reg_31_ ( .D(n447), .CK(clk), .Q(U1_C_31_) );
  DFF_X2 minm_reg_0_ ( .D(U5_Z_0), .CK(clk), .Q(minm[0]) );
  DFF_X2 minm_reg_11_ ( .D(U5_Z_11), .CK(clk), .Q(minm[11]) );
  DFF_X2 minm_reg_2_ ( .D(U5_Z_2), .CK(clk), .Q(minm[2]) );
  DFF_X2 in_cm_mac_reg_25_ ( .D(U6_Z_25), .CK(clk), .Q(U1_C_25_), .QN(n18) );
  DFF_X2 in_cm_mac_reg_27_ ( .D(U6_Z_27), .CK(clk), .Q(U1_C_27_), .QN(n12) );
  DFF_X2 in_cm_mac_reg_2_ ( .D(U6_Z_2), .CK(clk), .Q(U1_C_2_), .QN(n351) );
  DFF_X2 in_cm_mac_reg_0_ ( .D(U6_Z_0), .CK(clk), .Q(U1_C_0_), .QN(n513) );
  DFF_X2 in_cm_mac_reg_1_ ( .D(U6_Z_1), .CK(clk), .Q(U1_C_1_) );
  DFF_X2 in_cm_mac_reg_3_ ( .D(U6_Z_3), .CK(clk), .Q(U1_C_3_) );
  DFF_X2 in_cm_mac_reg_4_ ( .D(U6_Z_4), .CK(clk), .Q(U1_C_4_), .QN(n341) );
  DFF_X2 in_cm_mac_reg_6_ ( .D(U6_Z_6), .CK(clk), .Q(U1_C_6_) );
  DFF_X2 in_cm_mac_reg_7_ ( .D(U6_Z_7), .CK(clk), .Q(U1_C_7_) );
  DFF_X2 in_cm_mac_reg_8_ ( .D(U6_Z_8), .CK(clk), .Q(U1_C_8_), .QN(n678) );
  DFF_X2 in_cm_mac_reg_9_ ( .D(U6_Z_9), .CK(clk), .Q(U1_C_9_) );
  DFF_X2 in_cm_mac_reg_12_ ( .D(U6_Z_12), .CK(clk), .Q(U1_C_12_), .QN(n489) );
  DFF_X2 in_cm_mac_reg_10_ ( .D(U6_Z_10), .CK(clk), .Q(U1_C_10_), .QN(n498) );
  DFF_X2 in_cm_mac_reg_11_ ( .D(U6_Z_11), .CK(clk), .Q(U1_C_11_) );
  DFF_X2 in_cm_mac_reg_13_ ( .D(U6_Z_13), .CK(clk), .Q(U1_C_13_) );
  DFF_X2 in_cm_mac_reg_14_ ( .D(U6_Z_14), .CK(clk), .Q(U1_C_14_), .QN(n634) );
  DFF_X2 in_cm_mac_reg_15_ ( .D(U6_Z_15), .CK(clk), .Q(U1_C_15_) );
  DFF_X2 in_cm_mac_reg_16_ ( .D(U6_Z_16), .CK(clk), .Q(U1_C_16_) );
  DFF_X2 in_cm_mac_reg_18_ ( .D(U6_Z_18), .CK(clk), .Q(U1_C_18_) );
  DFF_X2 in_cm_mac_reg_20_ ( .D(U6_Z_20), .CK(clk), .Q(U1_C_20_) );
  DFF_X2 in_cm_mac_reg_22_ ( .D(U6_Z_22), .CK(clk), .Q(U1_C_22_) );
  DFF_X2 in_cm_mac_reg_24_ ( .D(U6_Z_24), .CK(clk), .Q(U1_C_24_) );
  DFF_X2 in_cm_mac_reg_28_ ( .D(U6_Z_28), .CK(clk), .Q(U1_C_28_) );
  DFF_X2 in_cm_mac_reg_5_ ( .D(U6_Z_5), .CK(clk), .Q(U1_C_5_), .QN(n280) );
  DFF_X2 in_cm_mac_reg_17_ ( .D(U6_Z_17), .CK(clk), .Q(U1_C_17_), .QN(n65) );
  DFF_X2 in_cm_mac_reg_19_ ( .D(U6_Z_19), .CK(clk), .Q(n609), .QN(n52) );
  DFF_X2 in_cm_mac_reg_21_ ( .D(U6_Z_21), .CK(clk), .Q(U1_C_21_), .QN(n41) );
  DFF_X2 in_cm_mac_reg_23_ ( .D(U6_Z_23), .CK(clk), .Q(U1_C_23_), .QN(n29) );
  DFF_X2 in_cm_mac_reg_29_ ( .D(U6_Z_29), .CK(clk), .Q(n1386), .QN(n4) );
  DFF_X2 minm_reg_5_ ( .D(U5_Z_5), .CK(clk), .Q(minm[5]) );
  DFF_X1 minm_reg_6_ ( .D(U5_Z_6), .CK(clk), .Q(minm[6]) );
  DFF_X1 minm_reg_1_ ( .D(U5_Z_1), .CK(clk), .Q(minm[1]) );
  DFF_X1 minm_reg_7_ ( .D(U5_Z_7), .CK(clk), .Q(minm[7]) );
  OAI22_X2 U8 ( .A1(n357), .A2(n1451), .B1(n1362), .B2(n1450), .ZN(n1370) );
  NAND2_X2 U10 ( .A1(n1005), .A2(n986), .ZN(n185) );
  NAND2_X2 U11 ( .A1(n183), .A2(n184), .ZN(n186) );
  NAND2_X2 U13 ( .A1(n185), .A2(n186), .ZN(n238) );
  INV_X4 U14 ( .A(n1005), .ZN(n183) );
  INV_X4 U15 ( .A(n986), .ZN(n184) );
  NAND2_X2 U16 ( .A1(n329), .A2(n504), .ZN(n189) );
  NAND2_X2 U17 ( .A1(n187), .A2(n188), .ZN(n190) );
  NAND2_X2 U18 ( .A1(n189), .A2(n190), .ZN(n254) );
  INV_X4 U19 ( .A(n329), .ZN(n187) );
  INV_X4 U20 ( .A(n504), .ZN(n188) );
  NAND2_X1 U21 ( .A1(n263), .A2(n192), .ZN(n193) );
  NAND2_X2 U22 ( .A1(n191), .A2(n1404), .ZN(n194) );
  NAND2_X2 U23 ( .A1(n193), .A2(n194), .ZN(n1399) );
  INV_X1 U24 ( .A(n263), .ZN(n191) );
  INV_X4 U25 ( .A(n1404), .ZN(n192) );
  OR2_X4 U26 ( .A1(n452), .A2(n1426), .ZN(n195) );
  OR2_X1 U27 ( .A1(n1283), .A2(n1282), .ZN(n196) );
  NAND2_X2 U28 ( .A1(n195), .A2(n196), .ZN(n288) );
  OAI22_X4 U38 ( .A1(n1273), .A2(n1272), .B1(n1271), .B2(n1270), .ZN(n1426) );
  INV_X1 U39 ( .A(n1427), .ZN(n1282) );
  INV_X4 U40 ( .A(n288), .ZN(n1430) );
  OAI21_X4 U46 ( .B1(n883), .B2(n1511), .A(n881), .ZN(n252) );
  NAND2_X4 U47 ( .A1(n456), .A2(n469), .ZN(n235) );
  NAND2_X2 U49 ( .A1(U1_C_3_), .A2(n529), .ZN(n551) );
  NOR2_X4 U50 ( .A1(n1491), .A2(n1490), .ZN(n1138) );
  INV_X4 U52 ( .A(n386), .ZN(n197) );
  INV_X8 U53 ( .A(in_z_mac[3]), .ZN(n1468) );
  NOR2_X4 U55 ( .A1(n1460), .A2(n1378), .ZN(n1383) );
  INV_X2 U56 ( .A(n1267), .ZN(n328) );
  NOR2_X2 U58 ( .A1(n1456), .A2(n1454), .ZN(n1369) );
  INV_X4 U59 ( .A(in_z_mac[7]), .ZN(n1572) );
  INV_X4 U61 ( .A(n440), .ZN(n455) );
  NAND2_X2 U62 ( .A1(n878), .A2(n876), .ZN(n881) );
  INV_X4 U63 ( .A(n386), .ZN(n457) );
  NOR2_X2 U64 ( .A1(n328), .A2(n1422), .ZN(n1265) );
  NOR2_X2 U65 ( .A1(n1452), .A2(n1357), .ZN(n1362) );
  OAI21_X2 U66 ( .B1(n592), .B2(n590), .A(n236), .ZN(n593) );
  INV_X4 U67 ( .A(n589), .ZN(n236) );
  NOR2_X2 U68 ( .A1(n1428), .A2(n1274), .ZN(n1283) );
  NOR2_X2 U69 ( .A1(n1521), .A2(n1522), .ZN(n1018) );
  NOR2_X2 U70 ( .A1(n1020), .A2(n1018), .ZN(n1487) );
  NAND2_X2 U71 ( .A1(n1409), .A2(n340), .ZN(n200) );
  NAND2_X2 U72 ( .A1(n198), .A2(n199), .ZN(n201) );
  NAND2_X2 U73 ( .A1(n200), .A2(n201), .ZN(n339) );
  INV_X4 U74 ( .A(n1409), .ZN(n198) );
  INV_X4 U75 ( .A(n340), .ZN(n199) );
  NAND2_X2 U76 ( .A1(n417), .A2(n584), .ZN(n204) );
  NAND2_X2 U77 ( .A1(n202), .A2(n203), .ZN(n205) );
  NAND2_X2 U78 ( .A1(n204), .A2(n205), .ZN(n589) );
  INV_X4 U79 ( .A(n417), .ZN(n202) );
  INV_X4 U80 ( .A(n584), .ZN(n203) );
  NOR2_X2 U81 ( .A1(n456), .A2(n581), .ZN(n206) );
  NOR2_X2 U82 ( .A1(n555), .A2(n235), .ZN(n207) );
  OR2_X2 U83 ( .A1(n206), .A2(n207), .ZN(n556) );
  INV_X4 U84 ( .A(n441), .ZN(n456) );
  INV_X2 U85 ( .A(n556), .ZN(n577) );
  NAND2_X2 U86 ( .A1(n389), .A2(n1154), .ZN(n211) );
  NAND2_X2 U87 ( .A1(n210), .A2(n1148), .ZN(n213) );
  NAND2_X2 U88 ( .A1(n211), .A2(n213), .ZN(n1141) );
  INV_X4 U89 ( .A(n389), .ZN(n210) );
  NOR2_X1 U90 ( .A1(n1149), .A2(n1148), .ZN(n1152) );
  INV_X1 U91 ( .A(n1456), .ZN(n297) );
  XNOR2_X2 U92 ( .A(n1016), .B(n402), .ZN(n1519) );
  OAI22_X1 U93 ( .A1(n1154), .A2(n1153), .B1(n1152), .B2(n1151), .ZN(n1162) );
  NOR2_X2 U94 ( .A1(n755), .A2(n752), .ZN(n1478) );
  AOI21_X2 U95 ( .B1(n816), .B2(n815), .A(n1574), .ZN(n710) );
  NAND2_X2 U96 ( .A1(n466), .A2(n1115), .ZN(n722) );
  OAI21_X2 U97 ( .B1(n1568), .B2(n1570), .A(n811), .ZN(n741) );
  OAI21_X2 U98 ( .B1(n733), .B2(n732), .A(n730), .ZN(n800) );
  NAND2_X2 U99 ( .A1(n464), .A2(n1125), .ZN(n815) );
  INV_X4 U100 ( .A(n321), .ZN(n322) );
  INV_X2 U101 ( .A(n292), .ZN(n293) );
  INV_X2 U102 ( .A(n1414), .ZN(n292) );
  XNOR2_X1 U103 ( .A(in_m_mac[14]), .B(n463), .ZN(n1063) );
  XNOR2_X1 U104 ( .A(in_m_mac[15]), .B(n463), .ZN(n1090) );
  XNOR2_X1 U105 ( .A(in_m_mac[13]), .B(n463), .ZN(n1056) );
  XNOR2_X1 U106 ( .A(in_m_mac[12]), .B(n463), .ZN(n1040) );
  XNOR2_X1 U107 ( .A(in_m_mac[11]), .B(n463), .ZN(n1012) );
  XNOR2_X1 U108 ( .A(in_m_mac[10]), .B(n463), .ZN(n981) );
  XNOR2_X1 U109 ( .A(in_m_mac[9]), .B(n463), .ZN(n950) );
  XNOR2_X1 U110 ( .A(in_m_mac[6]), .B(n463), .ZN(n830) );
  XNOR2_X1 U111 ( .A(in_m_mac[5]), .B(n463), .ZN(n817) );
  OAI21_X2 U112 ( .B1(n1571), .B2(n665), .A(n463), .ZN(n662) );
  XOR2_X1 U113 ( .A(n458), .B(n463), .Z(n717) );
  XOR2_X1 U114 ( .A(n463), .B(in_z_mac[8]), .Z(n1105) );
  NAND2_X1 U115 ( .A1(n459), .A2(n388), .ZN(n705) );
  AND2_X4 U116 ( .A1(n459), .A2(n386), .ZN(n214) );
  AND2_X4 U117 ( .A1(n585), .A2(n584), .ZN(n215) );
  INV_X1 U118 ( .A(n347), .ZN(n348) );
  INV_X2 U119 ( .A(n1420), .ZN(n347) );
  XOR2_X2 U120 ( .A(in_z_mac[14]), .B(in_z_mac[13]), .Z(n216) );
  AND2_X2 U121 ( .A1(n338), .A2(n337), .ZN(n218) );
  OAI22_X1 U122 ( .A1(n466), .A2(n985), .B1(n949), .B2(n722), .ZN(n983) );
  INV_X4 U123 ( .A(n228), .ZN(n1460) );
  INV_X4 U124 ( .A(n1403), .ZN(n263) );
  XNOR2_X2 U125 ( .A(n1385), .B(n300), .ZN(n219) );
  INV_X4 U126 ( .A(in_z_mac[5]), .ZN(n694) );
  XOR2_X2 U127 ( .A(in_z_mac[2]), .B(in_z_mac[3]), .Z(n220) );
  INV_X4 U128 ( .A(n458), .ZN(n459) );
  INV_X4 U129 ( .A(n444), .ZN(n464) );
  INV_X4 U130 ( .A(in_z_mac[0]), .ZN(n749) );
  INV_X4 U131 ( .A(n388), .ZN(n466) );
  XOR2_X1 U133 ( .A(in_z_mac[10]), .B(n463), .Z(n388) );
  INV_X4 U134 ( .A(n467), .ZN(n468) );
  XNOR2_X2 U135 ( .A(n1461), .B(n924), .ZN(n221) );
  NOR2_X2 U136 ( .A1(n823), .A2(n1235), .ZN(n222) );
  XNOR2_X2 U137 ( .A(n1445), .B(n371), .ZN(n223) );
  XNOR2_X2 U138 ( .A(n1292), .B(n960), .ZN(n224) );
  XNOR2_X2 U139 ( .A(n1306), .B(n993), .ZN(n225) );
  INV_X2 U140 ( .A(n1412), .ZN(n298) );
  AND2_X4 U141 ( .A1(n1122), .A2(n653), .ZN(n226) );
  OAI22_X2 U142 ( .A1(n1369), .A2(n1368), .B1(n1370), .B2(n1371), .ZN(n228) );
  INV_X2 U143 ( .A(n1252), .ZN(n1420) );
  INV_X4 U144 ( .A(n252), .ZN(n327) );
  INV_X2 U145 ( .A(n227), .ZN(n1155) );
  INV_X2 U146 ( .A(n1176), .ZN(n1502) );
  INV_X2 U147 ( .A(n1209), .ZN(n1509) );
  OAI22_X1 U148 ( .A1(n907), .A2(n905), .B1(n903), .B2(n902), .ZN(n969) );
  NAND2_X2 U149 ( .A1(n461), .A2(n749), .ZN(n240) );
  XNOR2_X1 U150 ( .A(in_m_mac[6]), .B(n461), .ZN(n575) );
  OAI22_X2 U151 ( .A1(n1237), .A2(n1238), .B1(n292), .B2(n1239), .ZN(n1252) );
  NAND2_X2 U152 ( .A1(n1497), .A2(n1156), .ZN(n227) );
  OAI22_X2 U153 ( .A1(n1383), .A2(n1382), .B1(n1458), .B2(n1384), .ZN(n229) );
  INV_X4 U154 ( .A(n229), .ZN(n1394) );
  NOR2_X1 U155 ( .A1(n439), .A2(n423), .ZN(U5_Z_14) );
  NOR2_X1 U156 ( .A1(n439), .A2(n258), .ZN(U5_Z_0) );
  XNOR2_X2 U157 ( .A(n1399), .B(n1401), .ZN(n423) );
  NOR2_X1 U158 ( .A1(n439), .A2(n243), .ZN(U5_Z_11) );
  NAND2_X1 U159 ( .A1(n1418), .A2(n1252), .ZN(n230) );
  INV_X2 U160 ( .A(n230), .ZN(n231) );
  OAI22_X2 U161 ( .A1(n1041), .A2(n1487), .B1(n1045), .B2(n1044), .ZN(n289) );
  OAI22_X2 U162 ( .A1(n1487), .A2(n1041), .B1(n1045), .B2(n1044), .ZN(n1491)
         );
  OAI22_X2 U163 ( .A1(n1264), .A2(n1265), .B1(n1266), .B2(n285), .ZN(n1284) );
  OAI22_X2 U164 ( .A1(n1174), .A2(n1499), .B1(n1176), .B2(n1175), .ZN(n1505)
         );
  OAI22_X1 U165 ( .A1(n214), .A2(n532), .B1(U1_C_2_), .B2(n533), .ZN(n546) );
  OAI22_X2 U166 ( .A1(n1208), .A2(n1507), .B1(n1508), .B2(n1209), .ZN(n1225)
         );
  XOR2_X2 U167 ( .A(n345), .B(n1572), .Z(n666) );
  INV_X2 U168 ( .A(n374), .ZN(n878) );
  INV_X1 U169 ( .A(n268), .ZN(n270) );
  INV_X1 U170 ( .A(n952), .ZN(n953) );
  XNOR2_X1 U171 ( .A(in_z_mac[5]), .B(n356), .ZN(n581) );
  INV_X4 U172 ( .A(n356), .ZN(n266) );
  XNOR2_X1 U173 ( .A(in_m_mac[2]), .B(in_z_mac[5]), .ZN(n753) );
  INV_X2 U174 ( .A(n935), .ZN(n681) );
  INV_X1 U175 ( .A(n310), .ZN(n232) );
  INV_X2 U176 ( .A(n553), .ZN(n310) );
  INV_X1 U177 ( .A(n566), .ZN(n233) );
  INV_X1 U178 ( .A(n344), .ZN(n345) );
  NAND2_X2 U179 ( .A1(n377), .A2(n378), .ZN(n441) );
  NOR2_X1 U180 ( .A1(n563), .A2(n341), .ZN(n564) );
  OAI22_X1 U181 ( .A1(n457), .A2(n684), .B1(n864), .B2(n364), .ZN(n935) );
  OAI22_X1 U182 ( .A1(n197), .A2(n1091), .B1(n1074), .B2(n362), .ZN(n1483) );
  OAI22_X1 U183 ( .A1(n1164), .A2(n362), .B1(n457), .B2(n1474), .ZN(n1477) );
  OAI22_X1 U184 ( .A1(n197), .A2(n1469), .B1(n1475), .B2(n362), .ZN(n1481) );
  OAI22_X1 U185 ( .A1(n457), .A2(n642), .B1(n640), .B2(n362), .ZN(n649) );
  NAND2_X2 U186 ( .A1(n456), .A2(n469), .ZN(n234) );
  XNOR2_X2 U187 ( .A(n857), .B(n856), .ZN(n241) );
  INV_X2 U188 ( .A(n749), .ZN(n321) );
  INV_X2 U189 ( .A(n437), .ZN(n313) );
  NAND2_X1 U190 ( .A1(n437), .A2(n422), .ZN(n315) );
  NAND2_X2 U191 ( .A1(n331), .A2(n332), .ZN(n237) );
  NAND2_X2 U192 ( .A1(n577), .A2(n578), .ZN(n331) );
  XNOR2_X2 U193 ( .A(n238), .B(n1003), .ZN(n1515) );
  OAI22_X1 U194 ( .A1(n962), .A2(n956), .B1(n954), .B2(n953), .ZN(n1003) );
  NAND2_X2 U195 ( .A1(n524), .A2(in_z_mac[3]), .ZN(n537) );
  INV_X4 U196 ( .A(n574), .ZN(n579) );
  OAI22_X2 U197 ( .A1(n197), .A2(n582), .B1(n559), .B2(n1473), .ZN(n574) );
  XNOR2_X2 U198 ( .A(n460), .B(n344), .ZN(n239) );
  INV_X2 U199 ( .A(n561), .ZN(n304) );
  NAND2_X2 U200 ( .A1(n461), .A2(n749), .ZN(n746) );
  INV_X4 U201 ( .A(in_z_mac[1]), .ZN(n543) );
  INV_X1 U202 ( .A(in_z_mac[1]), .ZN(n460) );
  NAND2_X1 U203 ( .A1(in_z_mac[5]), .A2(n459), .ZN(n308) );
  XOR2_X1 U204 ( .A(n694), .B(in_m_mac[3]), .Z(n754) );
  XOR2_X1 U205 ( .A(n694), .B(in_m_mac[5]), .Z(n716) );
  XOR2_X1 U206 ( .A(n694), .B(in_m_mac[6]), .Z(n695) );
  XOR2_X1 U207 ( .A(n694), .B(in_m_mac[9]), .Z(n492) );
  XOR2_X1 U208 ( .A(n694), .B(in_m_mac[10]), .Z(n474) );
  NAND2_X1 U209 ( .A1(n557), .A2(n234), .ZN(n558) );
  INV_X2 U210 ( .A(n828), .ZN(n819) );
  XOR2_X2 U211 ( .A(n356), .B(n1572), .Z(n596) );
  NAND2_X2 U212 ( .A1(in_z_mac[5]), .A2(n558), .ZN(n578) );
  XOR2_X1 U213 ( .A(in_m_mac[8]), .B(n1572), .Z(n831) );
  XNOR2_X1 U214 ( .A(in_m_mac[8]), .B(n463), .ZN(n901) );
  XOR2_X1 U215 ( .A(in_m_mac[8]), .B(n1573), .Z(n985) );
  XOR2_X1 U216 ( .A(in_m_mac[8]), .B(n1574), .Z(n1019) );
  XOR2_X1 U217 ( .A(in_m_mac[8]), .B(n1575), .Z(n1065) );
  XOR2_X1 U218 ( .A(n694), .B(in_m_mac[8]), .Z(n493) );
  NOR2_X2 U219 ( .A1(n459), .A2(n468), .ZN(n665) );
  NOR2_X2 U220 ( .A1(n208), .A2(n253), .ZN(n447) );
  XNOR2_X2 U221 ( .A(n241), .B(n759), .ZN(n902) );
  INV_X2 U222 ( .A(n759), .ZN(n858) );
  XNOR2_X1 U223 ( .A(in_z_mac[1]), .B(in_m_mac[1]), .ZN(n518) );
  INV_X4 U224 ( .A(n565), .ZN(n563) );
  INV_X1 U225 ( .A(n1571), .ZN(n246) );
  INV_X4 U226 ( .A(n643), .ZN(n1571) );
  NAND2_X2 U227 ( .A1(n468), .A2(n1105), .ZN(n643) );
  INV_X1 U228 ( .A(n538), .ZN(n251) );
  INV_X1 U229 ( .A(n541), .ZN(n538) );
  AOI21_X1 U230 ( .B1(n648), .B2(n647), .A(n645), .ZN(n715) );
  NOR2_X1 U231 ( .A1(n648), .A2(n647), .ZN(n497) );
  XOR2_X2 U232 ( .A(n1147), .B(n648), .Z(n381) );
  INV_X4 U233 ( .A(n832), .ZN(n883) );
  INV_X2 U234 ( .A(n439), .ZN(n253) );
  OAI21_X4 U235 ( .B1(n975), .B2(n1515), .A(n970), .ZN(n1521) );
  INV_X4 U236 ( .A(n254), .ZN(n1134) );
  INV_X2 U237 ( .A(n504), .ZN(n713) );
  NAND2_X1 U238 ( .A1(n441), .A2(n458), .ZN(n557) );
  XNOR2_X2 U239 ( .A(U1_C_7_), .B(n268), .ZN(n952) );
  OAI22_X1 U240 ( .A1(n946), .A2(n1462), .B1(n945), .B2(n455), .ZN(n912) );
  OAI22_X1 U241 ( .A1(n861), .A2(n1462), .B1(n946), .B2(n455), .ZN(n899) );
  OAI22_X1 U242 ( .A1(n1042), .A2(n1462), .B1(n1057), .B2(n455), .ZN(n1038) );
  OAI22_X1 U243 ( .A1(n977), .A2(n455), .B1(n945), .B2(n1462), .ZN(n630) );
  OAI22_X1 U244 ( .A1(n1017), .A2(n455), .B1(n977), .B2(n1462), .ZN(n613) );
  OAI22_X1 U245 ( .A1(n1042), .A2(n455), .B1(n1017), .B2(n1462), .ZN(n1278) );
  OAI22_X1 U246 ( .A1(n727), .A2(n455), .B1(n693), .B2(n1462), .ZN(n1107) );
  OAI22_X1 U247 ( .A1(n761), .A2(n455), .B1(n727), .B2(n1462), .ZN(n1143) );
  OAI22_X1 U248 ( .A1(n821), .A2(n455), .B1(n761), .B2(n1462), .ZN(n752) );
  OAI22_X1 U249 ( .A1(n831), .A2(n455), .B1(n821), .B2(n1462), .ZN(n478) );
  OAI22_X1 U250 ( .A1(n861), .A2(n455), .B1(n831), .B2(n1462), .ZN(n470) );
  AND2_X1 U251 ( .A1(n750), .A2(n1462), .ZN(n421) );
  NAND2_X1 U252 ( .A1(in_m_mac[2]), .A2(in_z_mac[1]), .ZN(n317) );
  INV_X4 U253 ( .A(in_z_mac[1]), .ZN(n387) );
  INV_X2 U254 ( .A(n1452), .ZN(n357) );
  NAND2_X2 U255 ( .A1(n267), .A2(n531), .ZN(n260) );
  NAND2_X1 U256 ( .A1(n267), .A2(n531), .ZN(n261) );
  INV_X1 U257 ( .A(n773), .ZN(n262) );
  INV_X1 U258 ( .A(n303), .ZN(n773) );
  NOR2_X1 U259 ( .A1(n352), .A2(n351), .ZN(n532) );
  NAND2_X2 U260 ( .A1(n457), .A2(n220), .ZN(n364) );
  NOR2_X1 U261 ( .A1(n516), .A2(n515), .ZN(n517) );
  AND2_X4 U262 ( .A1(n516), .A2(n515), .ZN(n349) );
  OAI22_X1 U263 ( .A1(n1136), .A2(n1135), .B1(n1134), .B2(n1133), .ZN(n1139)
         );
  INV_X1 U264 ( .A(n299), .ZN(n300) );
  INV_X1 U265 ( .A(n297), .ZN(n265) );
  INV_X4 U266 ( .A(n252), .ZN(n1516) );
  XNOR2_X2 U267 ( .A(n376), .B(in_z_mac[5]), .ZN(n469) );
  INV_X4 U268 ( .A(in_z_mac[4]), .ZN(n376) );
  INV_X4 U269 ( .A(n355), .ZN(n356) );
  INV_X1 U270 ( .A(n808), .ZN(n829) );
  INV_X2 U271 ( .A(n511), .ZN(n516) );
  XNOR2_X2 U272 ( .A(n519), .B(n214), .ZN(n267) );
  NOR2_X4 U273 ( .A1(n327), .A2(n1518), .ZN(n975) );
  XNOR2_X2 U274 ( .A(n460), .B(n344), .ZN(n544) );
  INV_X4 U275 ( .A(in_m_mac[3]), .ZN(n344) );
  OAI22_X1 U276 ( .A1(n468), .A2(n723), .B1(n692), .B2(n643), .ZN(n657) );
  OAI22_X1 U277 ( .A1(n468), .A2(n758), .B1(n723), .B2(n246), .ZN(n685) );
  OAI22_X1 U278 ( .A1(n468), .A2(n817), .B1(n758), .B2(n246), .ZN(n812) );
  OAI22_X1 U279 ( .A1(n641), .A2(n468), .B1(n643), .B2(n717), .ZN(n720) );
  XNOR2_X2 U280 ( .A(n892), .B(n868), .ZN(n1511) );
  OAI22_X1 U281 ( .A1(n854), .A2(n852), .B1(n851), .B2(n840), .ZN(n905) );
  OAI21_X2 U282 ( .B1(n549), .B2(n548), .A(n547), .ZN(n568) );
  INV_X4 U283 ( .A(n859), .ZN(n268) );
  INV_X1 U284 ( .A(n1487), .ZN(n271) );
  INV_X4 U285 ( .A(n271), .ZN(n272) );
  INV_X1 U286 ( .A(n878), .ZN(n273) );
  AND2_X1 U287 ( .A1(n579), .A2(n578), .ZN(n576) );
  INV_X1 U288 ( .A(n982), .ZN(n275) );
  INV_X1 U289 ( .A(n1005), .ZN(n982) );
  INV_X1 U290 ( .A(n234), .ZN(n276) );
  INV_X4 U291 ( .A(n276), .ZN(n277) );
  XNOR2_X1 U292 ( .A(n580), .B(n280), .ZN(n278) );
  INV_X4 U293 ( .A(n278), .ZN(n281) );
  XNOR2_X2 U294 ( .A(n1468), .B(n266), .ZN(n545) );
  INV_X1 U295 ( .A(n548), .ZN(n282) );
  INV_X4 U296 ( .A(n282), .ZN(n284) );
  OAI22_X2 U297 ( .A1(n347), .A2(n1418), .B1(n231), .B2(n1250), .ZN(n285) );
  INV_X1 U298 ( .A(n1521), .ZN(n286) );
  INV_X4 U299 ( .A(n286), .ZN(n287) );
  INV_X1 U300 ( .A(n1310), .ZN(n290) );
  INV_X1 U301 ( .A(n1349), .ZN(n291) );
  INV_X1 U302 ( .A(n1322), .ZN(n295) );
  INV_X1 U303 ( .A(n263), .ZN(n296) );
  INV_X2 U304 ( .A(n1444), .ZN(n370) );
  INV_X2 U305 ( .A(n1428), .ZN(n452) );
  INV_X1 U306 ( .A(n1394), .ZN(n299) );
  XNOR2_X2 U307 ( .A(in_z_mac[7]), .B(in_z_mac[8]), .ZN(n614) );
  INV_X4 U308 ( .A(n764), .ZN(n768) );
  INV_X2 U309 ( .A(n240), .ZN(n301) );
  INV_X4 U310 ( .A(n301), .ZN(n302) );
  XNOR2_X2 U311 ( .A(n808), .B(n825), .ZN(n325) );
  XNOR2_X2 U312 ( .A(n688), .B(n418), .ZN(n303) );
  XOR2_X2 U313 ( .A(n409), .B(n937), .Z(n986) );
  NAND2_X1 U314 ( .A1(n237), .A2(n574), .ZN(n305) );
  NAND2_X2 U315 ( .A1(n304), .A2(n579), .ZN(n306) );
  NAND2_X2 U316 ( .A1(n305), .A2(n306), .ZN(n326) );
  NAND2_X1 U317 ( .A1(n694), .A2(n458), .ZN(n307) );
  NAND2_X2 U318 ( .A1(n307), .A2(n308), .ZN(n555) );
  NAND2_X1 U319 ( .A1(n551), .A2(n553), .ZN(n311) );
  NAND2_X2 U320 ( .A1(n309), .A2(n310), .ZN(n312) );
  NAND2_X2 U321 ( .A1(n311), .A2(n312), .ZN(n350) );
  INV_X1 U322 ( .A(n551), .ZN(n309) );
  NAND2_X2 U323 ( .A1(n313), .A2(n314), .ZN(n316) );
  NAND2_X2 U324 ( .A1(n315), .A2(n316), .ZN(n553) );
  INV_X1 U325 ( .A(n422), .ZN(n314) );
  OAI22_X2 U326 ( .A1(n309), .A2(n554), .B1(n232), .B2(n552), .ZN(n588) );
  INV_X2 U327 ( .A(n833), .ZN(n854) );
  XNOR2_X2 U328 ( .A(in_m_mac[5]), .B(n461), .ZN(n560) );
  XNOR2_X2 U329 ( .A(n867), .B(U1_C_6_), .ZN(n436) );
  AND2_X4 U330 ( .A1(n867), .A2(U1_C_6_), .ZN(n866) );
  OAI22_X2 U331 ( .A1(n459), .A2(n240), .B1(n518), .B2(n322), .ZN(n510) );
  NAND2_X2 U332 ( .A1(n585), .A2(n281), .ZN(n359) );
  INV_X2 U333 ( .A(n326), .ZN(n585) );
  NAND2_X2 U334 ( .A1(n387), .A2(n319), .ZN(n318) );
  NAND2_X2 U335 ( .A1(n317), .A2(n318), .ZN(n528) );
  INV_X1 U337 ( .A(in_m_mac[2]), .ZN(n319) );
  INV_X2 U338 ( .A(n319), .ZN(n320) );
  NAND2_X1 U339 ( .A1(n586), .A2(n326), .ZN(n587) );
  NAND2_X1 U340 ( .A1(n326), .A2(n278), .ZN(n360) );
  INV_X1 U341 ( .A(n789), .ZN(n323) );
  INV_X4 U342 ( .A(n323), .ZN(n324) );
  XNOR2_X2 U343 ( .A(n833), .B(n448), .ZN(n583) );
  XNOR2_X2 U344 ( .A(n325), .B(n828), .ZN(n788) );
  XOR2_X1 U345 ( .A(in_m_mac[4]), .B(n1574), .Z(n894) );
  XOR2_X1 U346 ( .A(in_m_mac[4]), .B(n1575), .Z(n984) );
  INV_X2 U347 ( .A(n1511), .ZN(n1512) );
  NAND2_X1 U348 ( .A1(U1_C_7_), .A2(n270), .ZN(n762) );
  NAND3_X2 U349 ( .A1(U1_C_7_), .A2(n768), .A3(n270), .ZN(n915) );
  NOR2_X4 U350 ( .A1(n1444), .A2(n1333), .ZN(n1334) );
  NOR2_X4 U351 ( .A1(n1412), .A2(n1410), .ZN(n1223) );
  INV_X4 U352 ( .A(n1284), .ZN(n1428) );
  OAI22_X1 U353 ( .A1(n834), .A2(n322), .B1(n818), .B2(n302), .ZN(n639) );
  OAI22_X1 U354 ( .A1(n897), .A2(n322), .B1(n834), .B2(n302), .ZN(n1464) );
  OAI21_X2 U355 ( .B1(n1138), .B2(n1492), .A(n1137), .ZN(n1497) );
  XOR2_X1 U356 ( .A(n694), .B(in_m_mac[7]), .Z(n494) );
  XOR2_X1 U357 ( .A(in_m_mac[7]), .B(n1572), .Z(n821) );
  XNOR2_X1 U358 ( .A(in_m_mac[7]), .B(n463), .ZN(n874) );
  XOR2_X1 U359 ( .A(in_m_mac[7]), .B(n1573), .Z(n949) );
  XOR2_X1 U360 ( .A(n1573), .B(n459), .Z(n726) );
  XOR2_X1 U361 ( .A(n1574), .B(n459), .Z(n814) );
  XOR2_X1 U362 ( .A(n1575), .B(n459), .Z(n873) );
  NAND2_X1 U363 ( .A1(n321), .A2(n459), .ZN(n514) );
  NAND2_X1 U364 ( .A1(n459), .A2(n216), .ZN(n633) );
  AND2_X4 U365 ( .A1(n441), .A2(n459), .ZN(n422) );
  INV_X1 U366 ( .A(n285), .ZN(n1424) );
  XOR2_X1 U367 ( .A(n595), .B(n324), .Z(n598) );
  XNOR2_X2 U368 ( .A(n712), .B(n636), .ZN(n329) );
  OAI22_X2 U369 ( .A1(n456), .A2(n753), .B1(n581), .B2(n235), .ZN(n840) );
  NAND2_X2 U370 ( .A1(n556), .A2(n330), .ZN(n332) );
  NAND2_X2 U371 ( .A1(n331), .A2(n332), .ZN(n561) );
  INV_X2 U372 ( .A(n578), .ZN(n330) );
  BUF_X4 U373 ( .A(n1497), .Z(n333) );
  NOR2_X2 U374 ( .A1(n263), .A2(n1400), .ZN(n1402) );
  NOR2_X2 U375 ( .A1(n1439), .A2(n1316), .ZN(n1321) );
  XNOR2_X1 U376 ( .A(in_m_mac[7]), .B(n461), .ZN(n591) );
  XNOR2_X1 U377 ( .A(in_m_mac[8]), .B(n461), .ZN(n615) );
  XNOR2_X1 U378 ( .A(in_m_mac[10]), .B(n461), .ZN(n697) );
  XNOR2_X1 U379 ( .A(in_m_mac[12]), .B(n461), .ZN(n747) );
  XNOR2_X1 U380 ( .A(in_m_mac[14]), .B(n461), .ZN(n834) );
  XNOR2_X1 U381 ( .A(in_m_mac[15]), .B(n461), .ZN(n897) );
  XNOR2_X1 U382 ( .A(in_m_mac[13]), .B(n461), .ZN(n818) );
  XNOR2_X1 U383 ( .A(in_m_mac[11]), .B(n461), .ZN(n748) );
  XNOR2_X1 U384 ( .A(in_m_mac[9]), .B(n461), .ZN(n661) );
  NAND2_X1 U385 ( .A1(n572), .A2(n571), .ZN(n334) );
  INV_X2 U386 ( .A(n568), .ZN(n566) );
  OAI22_X1 U387 ( .A1(n456), .A2(n754), .B1(n753), .B2(n235), .ZN(n856) );
  NAND2_X1 U388 ( .A1(n350), .A2(n554), .ZN(n337) );
  NAND2_X2 U389 ( .A1(n335), .A2(n336), .ZN(n338) );
  INV_X2 U390 ( .A(n350), .ZN(n335) );
  INV_X1 U391 ( .A(n554), .ZN(n336) );
  OAI22_X1 U392 ( .A1(n197), .A2(n559), .B1(n362), .B2(n545), .ZN(n554) );
  INV_X4 U393 ( .A(n339), .ZN(n439) );
  XOR2_X2 U394 ( .A(U1_C_31_), .B(n1408), .Z(n340) );
  OAI22_X1 U395 ( .A1(n457), .A2(n640), .B1(n1469), .B2(n362), .ZN(n1218) );
  OAI22_X1 U396 ( .A1(n457), .A2(n1475), .B1(n1474), .B2(n1473), .ZN(n1482) );
  OAI22_X1 U397 ( .A1(n197), .A2(n1164), .B1(n1091), .B2(n362), .ZN(n1168) );
  INV_X2 U398 ( .A(n537), .ZN(n542) );
  NOR2_X1 U399 ( .A1(n538), .A2(n537), .ZN(n539) );
  OAI22_X1 U400 ( .A1(n457), .A2(n1074), .B1(n686), .B2(n1473), .ZN(n504) );
  OAI22_X1 U401 ( .A1(n457), .A2(n860), .B1(n582), .B2(n364), .ZN(n852) );
  OAI21_X4 U402 ( .B1(n527), .B2(n1473), .A(n526), .ZN(n541) );
  NAND2_X2 U403 ( .A1(n197), .A2(n220), .ZN(n1473) );
  OAI22_X2 U404 ( .A1(n239), .A2(n322), .B1(n746), .B2(n528), .ZN(n529) );
  NAND2_X1 U405 ( .A1(n565), .A2(U1_C_4_), .ZN(n342) );
  NAND2_X2 U406 ( .A1(n563), .A2(n341), .ZN(n343) );
  NAND2_X2 U407 ( .A1(n342), .A2(n343), .ZN(n437) );
  INV_X4 U408 ( .A(n298), .ZN(n346) );
  XNOR2_X1 U409 ( .A(n459), .B(in_z_mac[3]), .ZN(n527) );
  OAI22_X1 U410 ( .A1(n514), .A2(n513), .B1(n512), .B2(n387), .ZN(n515) );
  NOR2_X2 U411 ( .A1(n546), .A2(n260), .ZN(n549) );
  NAND2_X1 U412 ( .A1(n533), .A2(U1_C_2_), .ZN(n353) );
  NAND2_X2 U413 ( .A1(n351), .A2(n352), .ZN(n354) );
  NAND2_X2 U414 ( .A1(n353), .A2(n354), .ZN(n519) );
  INV_X2 U415 ( .A(n533), .ZN(n352) );
  INV_X1 U416 ( .A(in_m_mac[1]), .ZN(n355) );
  INV_X2 U417 ( .A(n357), .ZN(n358) );
  NAND2_X2 U418 ( .A1(n359), .A2(n360), .ZN(n417) );
  NAND2_X2 U419 ( .A1(n457), .A2(n220), .ZN(n362) );
  INV_X1 U420 ( .A(n375), .ZN(n365) );
  INV_X1 U422 ( .A(n556), .ZN(n366) );
  INV_X4 U423 ( .A(n370), .ZN(n371) );
  INV_X1 U424 ( .A(n1509), .ZN(n372) );
  INV_X4 U425 ( .A(n372), .ZN(n373) );
  NAND2_X2 U426 ( .A1(n1516), .A2(n1518), .ZN(n970) );
  NAND2_X2 U427 ( .A1(n793), .A2(n805), .ZN(n374) );
  OAI21_X4 U428 ( .B1(n789), .B2(n791), .A(n788), .ZN(n793) );
  NOR2_X1 U429 ( .A1(n625), .A2(n624), .ZN(n1167) );
  NAND2_X2 U430 ( .A1(n1468), .A2(in_z_mac[4]), .ZN(n377) );
  INV_X1 U431 ( .A(n1182), .ZN(n375) );
  XOR2_X1 U432 ( .A(n1468), .B(in_m_mac[5]), .Z(n864) );
  XOR2_X1 U433 ( .A(n1468), .B(in_m_mac[4]), .Z(n860) );
  INV_X2 U434 ( .A(n1177), .ZN(n1181) );
  NOR2_X2 U435 ( .A1(n806), .A2(n807), .ZN(n1470) );
  AND2_X1 U436 ( .A1(n780), .A2(n778), .ZN(n1476) );
  XNOR2_X2 U437 ( .A(n381), .B(n647), .ZN(n1157) );
  INV_X4 U438 ( .A(n1135), .ZN(n419) );
  AOI21_X2 U439 ( .B1(n721), .B2(n722), .A(n1573), .ZN(n658) );
  XOR2_X2 U442 ( .A(n782), .B(n781), .Z(n382) );
  AND2_X4 U443 ( .A1(n459), .A2(n467), .ZN(n428) );
  NAND2_X2 U444 ( .A1(n465), .A2(n1123), .ZN(n361) );
  INV_X4 U445 ( .A(in_z_mac[11]), .ZN(n1573) );
  NAND2_X2 U446 ( .A1(in_z_mac[3]), .A2(n376), .ZN(n378) );
  AND2_X4 U447 ( .A1(n1180), .A2(n1181), .ZN(n1178) );
  OAI21_X2 U448 ( .B1(n710), .B2(n812), .A(n711), .ZN(n811) );
  XNOR2_X1 U449 ( .A(n935), .B(n934), .ZN(n409) );
  XOR2_X2 U450 ( .A(n379), .B(n1203), .Z(n1196) );
  XOR2_X2 U451 ( .A(n1204), .B(n380), .Z(n379) );
  XOR2_X1 U452 ( .A(n1460), .B(n413), .Z(n242) );
  XNOR2_X1 U453 ( .A(n708), .B(n677), .ZN(n676) );
  INV_X1 U454 ( .A(n1139), .ZN(n398) );
  NOR2_X1 U455 ( .A1(n657), .A2(n658), .ZN(n1484) );
  AND2_X4 U456 ( .A1(n687), .A2(n685), .ZN(n484) );
  AOI21_X1 U458 ( .B1(n770), .B2(n222), .A(n767), .ZN(n795) );
  NOR2_X1 U459 ( .A1(n770), .A2(n222), .ZN(n1236) );
  NAND2_X1 U460 ( .A1(n431), .A2(n736), .ZN(n1217) );
  INV_X1 U461 ( .A(n677), .ZN(n1526) );
  AOI21_X1 U462 ( .B1(n842), .B2(n843), .A(n841), .ZN(n885) );
  NOR2_X1 U463 ( .A1(n843), .A2(n842), .ZN(n1262) );
  INV_X2 U464 ( .A(n545), .ZN(n525) );
  OR2_X4 U465 ( .A1(n421), .A2(n1572), .ZN(n857) );
  XNOR2_X2 U467 ( .A(n809), .B(n424), .ZN(n380) );
  XNOR2_X1 U468 ( .A(n625), .B(n624), .ZN(n427) );
  XNOR2_X2 U469 ( .A(n382), .B(n783), .ZN(n1006) );
  AOI21_X1 U470 ( .B1(n869), .B2(n361), .A(n1575), .ZN(n807) );
  NOR2_X1 U471 ( .A1(n776), .A2(n824), .ZN(n1235) );
  INV_X1 U472 ( .A(n900), .ZN(n1534) );
  OAI21_X1 U473 ( .B1(n1563), .B2(n900), .A(n947), .ZN(n886) );
  XNOR2_X1 U474 ( .A(n1508), .B(n1507), .ZN(n1510) );
  XOR2_X1 U475 ( .A(n1506), .B(n365), .Z(n264) );
  XNOR2_X1 U476 ( .A(n1504), .B(n1503), .ZN(n1506) );
  XOR2_X1 U477 ( .A(n1500), .B(n1499), .Z(n1501) );
  XOR2_X1 U478 ( .A(n383), .B(n1522), .Z(n209) );
  XNOR2_X1 U479 ( .A(n287), .B(n1520), .ZN(n383) );
  XNOR2_X1 U480 ( .A(n1490), .B(n1494), .ZN(n279) );
  XOR2_X1 U481 ( .A(n1493), .B(n1492), .Z(n1494) );
  XOR2_X1 U482 ( .A(n384), .B(n1514), .Z(n217) );
  XNOR2_X1 U483 ( .A(n273), .B(n1512), .ZN(n384) );
  XNOR2_X1 U484 ( .A(n1515), .B(n451), .ZN(n1517) );
  XOR2_X1 U485 ( .A(n1518), .B(n1517), .Z(n212) );
  XNOR2_X1 U487 ( .A(n385), .B(n592), .ZN(n573) );
  XOR2_X1 U488 ( .A(n588), .B(n589), .Z(n385) );
  XNOR2_X1 U489 ( .A(n569), .B(n218), .ZN(n435) );
  XOR2_X1 U490 ( .A(n435), .B(n233), .Z(n550) );
  XOR2_X1 U491 ( .A(n534), .B(n546), .Z(n535) );
  XNOR2_X2 U492 ( .A(in_z_mac[2]), .B(n543), .ZN(n386) );
  XNOR2_X1 U493 ( .A(in_m_mac[13]), .B(in_z_mac[5]), .ZN(n644) );
  INV_X4 U494 ( .A(n216), .ZN(n465) );
  XNOR2_X1 U496 ( .A(in_m_mac[14]), .B(in_z_mac[5]), .ZN(n619) );
  XNOR2_X2 U497 ( .A(n1150), .B(n1149), .ZN(n389) );
  XNOR2_X2 U498 ( .A(n390), .B(n1210), .ZN(n1507) );
  XNOR2_X2 U499 ( .A(n1212), .B(n1216), .ZN(n390) );
  XNOR2_X2 U500 ( .A(n391), .B(n1194), .ZN(n1504) );
  XNOR2_X2 U501 ( .A(n1196), .B(n1200), .ZN(n391) );
  XNOR2_X2 U502 ( .A(n392), .B(n1158), .ZN(n1496) );
  XNOR2_X2 U503 ( .A(n1159), .B(n1163), .ZN(n392) );
  XNOR2_X2 U504 ( .A(n393), .B(n1181), .ZN(n1499) );
  XNOR2_X2 U505 ( .A(n1180), .B(n1179), .ZN(n393) );
  XOR2_X2 U506 ( .A(n794), .B(n394), .Z(n1242) );
  XNOR2_X2 U507 ( .A(n1529), .B(n1551), .ZN(n394) );
  XNOR2_X2 U508 ( .A(n1226), .B(n395), .ZN(n1411) );
  XNOR2_X2 U509 ( .A(n414), .B(n1227), .ZN(n395) );
  XNOR2_X2 U510 ( .A(n396), .B(n1241), .ZN(n1415) );
  XNOR2_X2 U511 ( .A(n1242), .B(n1240), .ZN(n396) );
  XNOR2_X2 U512 ( .A(n1443), .B(n1442), .ZN(n1445) );
  OR2_X1 U514 ( .A1(n845), .A2(n397), .ZN(n1253) );
  AND2_X4 U515 ( .A1(n844), .A2(n1529), .ZN(n397) );
  AOI21_X2 U517 ( .B1(n846), .B2(n1551), .A(n794), .ZN(n845) );
  XNOR2_X2 U518 ( .A(n902), .B(n895), .ZN(n868) );
  XNOR2_X2 U519 ( .A(n399), .B(n398), .ZN(n1492) );
  XNOR2_X2 U520 ( .A(n1142), .B(n1141), .ZN(n399) );
  XNOR2_X2 U521 ( .A(n400), .B(n738), .ZN(n1045) );
  XNOR2_X2 U522 ( .A(n737), .B(n735), .ZN(n400) );
  XNOR2_X2 U523 ( .A(n401), .B(n1119), .ZN(n1153) );
  XNOR2_X2 U524 ( .A(n1107), .B(n654), .ZN(n401) );
  XNOR2_X2 U525 ( .A(n303), .B(n1015), .ZN(n402) );
  XNOR2_X2 U526 ( .A(n403), .B(n704), .ZN(n739) );
  XNOR2_X2 U527 ( .A(n696), .B(n1569), .ZN(n403) );
  OAI22_X1 U528 ( .A1(n636), .A2(n504), .B1(n503), .B2(n712), .ZN(n625) );
  AND2_X1 U529 ( .A1(n1142), .A2(n398), .ZN(n1140) );
  XNOR2_X2 U532 ( .A(n404), .B(n479), .ZN(n699) );
  XNOR2_X2 U533 ( .A(n478), .B(n784), .ZN(n404) );
  XNOR2_X2 U536 ( .A(n405), .B(n674), .ZN(n1180) );
  XNOR2_X2 U537 ( .A(n673), .B(n1189), .ZN(n405) );
  XNOR2_X2 U538 ( .A(n1172), .B(n406), .ZN(n1159) );
  XNOR2_X2 U539 ( .A(n1525), .B(n1524), .ZN(n406) );
  XNOR2_X2 U540 ( .A(n734), .B(n407), .ZN(n1212) );
  XNOR2_X2 U541 ( .A(n736), .B(n431), .ZN(n407) );
  XNOR2_X2 U543 ( .A(n1483), .B(n408), .ZN(n1150) );
  XNOR2_X2 U544 ( .A(n657), .B(n658), .ZN(n408) );
  AOI21_X1 U545 ( .B1(n657), .B2(n658), .A(n1564), .ZN(n648) );
  AOI21_X1 U546 ( .B1(n755), .B2(n752), .A(n1559), .ZN(n809) );
  AND2_X1 U547 ( .A1(n496), .A2(n654), .ZN(n495) );
  AND2_X1 U548 ( .A1(n865), .A2(n863), .ZN(n1467) );
  XNOR2_X2 U549 ( .A(n410), .B(n806), .ZN(n733) );
  XNOR2_X2 U550 ( .A(n1481), .B(n807), .ZN(n410) );
  AOI21_X1 U551 ( .B1(n732), .B2(n733), .A(n1527), .ZN(n770) );
  AOI21_X2 U552 ( .B1(n1530), .B2(n849), .A(n890), .ZN(n842) );
  AOI21_X2 U553 ( .B1(n891), .B2(n1548), .A(n848), .ZN(n890) );
  XOR2_X2 U554 ( .A(n863), .B(n411), .Z(n796) );
  XNOR2_X2 U557 ( .A(n1472), .B(n865), .ZN(n411) );
  AOI21_X2 U558 ( .B1(n912), .B2(n909), .A(n1557), .ZN(n888) );
  OAI21_X2 U559 ( .B1(n909), .B2(n912), .A(n911), .ZN(n942) );
  AOI21_X1 U560 ( .B1(n804), .B2(n801), .A(n1566), .ZN(n798) );
  OAI21_X1 U561 ( .B1(n801), .B2(n804), .A(n803), .ZN(n871) );
  AOI21_X1 U563 ( .B1(n806), .B2(n807), .A(n1552), .ZN(n799) );
  XOR2_X2 U565 ( .A(n841), .B(n412), .Z(n1256) );
  XOR2_X2 U566 ( .A(n842), .B(n843), .Z(n412) );
  XOR2_X2 U567 ( .A(n1459), .B(n1458), .Z(n413) );
  OAI21_X1 U568 ( .B1(n431), .B2(n736), .A(n734), .ZN(n771) );
  OAI21_X1 U569 ( .B1(n766), .B2(n765), .A(n763), .ZN(n850) );
  OAI21_X1 U570 ( .B1(n1526), .B2(n708), .A(n675), .ZN(n707) );
  XNOR2_X2 U571 ( .A(n767), .B(n415), .ZN(n414) );
  XNOR2_X2 U572 ( .A(n222), .B(n770), .ZN(n415) );
  AOI21_X2 U573 ( .B1(n974), .B2(n971), .A(n1556), .ZN(n921) );
  OAI21_X2 U574 ( .B1(n971), .B2(n974), .A(n973), .ZN(n1009) );
  AOI21_X2 U575 ( .B1(n1001), .B2(n998), .A(n1555), .ZN(n989) );
  OAI21_X2 U576 ( .B1(n998), .B2(n1001), .A(n1000), .ZN(n1058) );
  OAI21_X2 U577 ( .B1(n997), .B2(n1539), .A(n959), .ZN(n996) );
  OAI21_X2 U578 ( .B1(n925), .B2(n1536), .A(n923), .ZN(n963) );
  OAI21_X2 U579 ( .B1(n1561), .B2(n1033), .A(n1064), .ZN(n1027) );
  OAI21_X2 U580 ( .B1(n1032), .B2(n1547), .A(n1034), .ZN(n1064) );
  OAI21_X2 U581 ( .B1(n1086), .B2(n1560), .A(n1101), .ZN(n1078) );
  OAI21_X2 U582 ( .B1(n1102), .B2(n1546), .A(n1087), .ZN(n1101) );
  XNOR2_X2 U583 ( .A(n416), .B(n951), .ZN(n907) );
  XNOR2_X2 U585 ( .A(n952), .B(n962), .ZN(n416) );
  XNOR2_X2 U586 ( .A(n743), .B(n742), .ZN(n418) );
  XNOR2_X2 U587 ( .A(n420), .B(n419), .ZN(n737) );
  XNOR2_X2 U588 ( .A(n1134), .B(n1132), .ZN(n420) );
  AND2_X1 U591 ( .A1(n1136), .A2(n1135), .ZN(n1133) );
  XNOR2_X2 U592 ( .A(n740), .B(n741), .ZN(n424) );
  AOI21_X2 U593 ( .B1(n699), .B2(n701), .A(n702), .ZN(n777) );
  XNOR2_X2 U594 ( .A(n425), .B(n1183), .ZN(n677) );
  XNOR2_X2 U597 ( .A(n1184), .B(n1185), .ZN(n425) );
  XOR2_X2 U598 ( .A(n426), .B(n1130), .Z(n728) );
  XNOR2_X2 U599 ( .A(n1126), .B(n1128), .ZN(n426) );
  XNOR2_X2 U600 ( .A(n427), .B(n622), .ZN(n1142) );
  OAI21_X2 U601 ( .B1(n215), .B2(n281), .A(n587), .ZN(n786) );
  AOI21_X1 U602 ( .B1(n625), .B2(n624), .A(n622), .ZN(n689) );
  AND2_X1 U603 ( .A1(n720), .A2(n782), .ZN(n719) );
  XNOR2_X2 U605 ( .A(n1398), .B(n1397), .ZN(n1385) );
  AND2_X1 U606 ( .A1(n459), .A2(n440), .ZN(n429) );
  AOI21_X2 U607 ( .B1(n790), .B2(n1261), .A(n908), .ZN(n843) );
  AOI21_X2 U608 ( .B1(n1532), .B2(n1538), .A(n792), .ZN(n908) );
  OAI21_X1 U609 ( .B1(n809), .B2(n740), .A(n810), .ZN(n732) );
  OAI21_X1 U610 ( .B1(n1528), .B2(n1558), .A(n741), .ZN(n810) );
  AOI21_X1 U611 ( .B1(n855), .B2(n1535), .A(n1531), .ZN(n891) );
  OAI21_X2 U613 ( .B1(n1535), .B2(n855), .A(n446), .ZN(n896) );
  XOR2_X2 U614 ( .A(n430), .B(n699), .Z(n1195) );
  XNOR2_X2 U615 ( .A(n1190), .B(n702), .ZN(n430) );
  AOI21_X2 U617 ( .B1(n838), .B2(n836), .A(n1537), .ZN(n884) );
  OAI21_X2 U618 ( .B1(n836), .B2(n838), .A(n839), .ZN(n931) );
  AOI21_X1 U619 ( .B1(n197), .B2(n1473), .A(n642), .ZN(n1463) );
  AOI21_X2 U622 ( .B1(n880), .B2(n879), .A(n877), .ZN(n968) );
  XNOR2_X2 U623 ( .A(n824), .B(n774), .ZN(n431) );
  AOI21_X1 U624 ( .B1(n824), .B2(n776), .A(n775), .ZN(n823) );
  AOI21_X2 U625 ( .B1(n886), .B2(n1275), .A(n941), .ZN(n1523) );
  AOI21_X2 U626 ( .B1(n1533), .B2(n889), .A(n888), .ZN(n941) );
  OAI21_X2 U628 ( .B1(n965), .B2(n966), .A(n967), .ZN(n1013) );
  OAI21_X2 U629 ( .B1(n927), .B2(n930), .A(n929), .ZN(n979) );
  OAI21_X2 U632 ( .B1(n1534), .B2(n948), .A(n914), .ZN(n947) );
  OR2_X1 U633 ( .A1(n432), .A2(n897), .ZN(n626) );
  AND2_X4 U634 ( .A1(n302), .A2(n322), .ZN(n432) );
  AOI21_X2 U635 ( .B1(n958), .B2(n957), .A(n955), .ZN(n1035) );
  OR2_X1 U637 ( .A1(n433), .A2(n1057), .ZN(n1547) );
  AND2_X4 U639 ( .A1(n455), .A2(n1462), .ZN(n433) );
  OAI21_X2 U640 ( .B1(n1550), .B2(n989), .A(n1542), .ZN(n1028) );
  AOI21_X2 U641 ( .B1(n989), .B2(n1550), .A(n991), .ZN(n1054) );
  OAI21_X2 U642 ( .B1(n995), .B2(n994), .A(n992), .ZN(n1029) );
  AOI21_X2 U643 ( .B1(n1049), .B2(n1048), .A(n1046), .ZN(n1082) );
  OAI21_X2 U644 ( .B1(n1028), .B2(n1027), .A(n1025), .ZN(n1050) );
  OAI21_X2 U645 ( .B1(n1022), .B2(n1023), .A(n1024), .ZN(n1068) );
  AOI21_X1 U646 ( .B1(n722), .B2(n466), .A(n1112), .ZN(n1096) );
  AOI21_X2 U647 ( .B1(n1095), .B2(n1553), .A(n1096), .ZN(n1111) );
  OAI21_X2 U648 ( .B1(n1078), .B2(n1081), .A(n1080), .ZN(n1098) );
  XNOR2_X2 U649 ( .A(n454), .B(n1501), .ZN(n269) );
  OR2_X1 U650 ( .A1(n434), .A2(n1124), .ZN(n655) );
  AND2_X4 U651 ( .A1(n815), .A2(n464), .ZN(n434) );
  XNOR2_X2 U652 ( .A(n436), .B(n429), .ZN(n825) );
  XNOR2_X2 U655 ( .A(n438), .B(n706), .ZN(n1132) );
  XNOR2_X2 U656 ( .A(n705), .B(U1_C_10_), .ZN(n438) );
  OAI21_X2 U657 ( .B1(U1_C_3_), .B2(n529), .A(n551), .ZN(n536) );
  INV_X4 U658 ( .A(in_m_mac[0]), .ZN(n458) );
  INV_X8 U659 ( .A(n462), .ZN(n463) );
  INV_X4 U664 ( .A(in_z_mac[9]), .ZN(n462) );
  XOR2_X2 U665 ( .A(in_z_mac[6]), .B(in_z_mac[5]), .Z(n440) );
  OAI21_X1 U666 ( .B1(U1_C_1_), .B2(n510), .A(n520), .ZN(n511) );
  INV_X4 U667 ( .A(n614), .ZN(n467) );
  XNOR2_X2 U668 ( .A(n442), .B(n428), .ZN(n918) );
  XNOR2_X2 U670 ( .A(n745), .B(U1_C_8_), .ZN(n442) );
  XNOR2_X2 U672 ( .A(n443), .B(n506), .ZN(n1147) );
  XNOR2_X2 U673 ( .A(n505), .B(U1_C_12_), .ZN(n443) );
  OAI21_X2 U675 ( .B1(U1_C_11_), .B2(n507), .A(n1144), .ZN(n622) );
  XNOR2_X2 U676 ( .A(in_z_mac[12]), .B(n1573), .ZN(n444) );
  XNOR2_X2 U679 ( .A(n445), .B(n635), .ZN(n1190) );
  XNOR2_X2 U680 ( .A(n633), .B(U1_C_14_), .ZN(n445) );
  INV_X4 U682 ( .A(in_z_mac[13]), .ZN(n1574) );
  INV_X4 U683 ( .A(in_z_mac[15]), .ZN(n1575) );
  AOI21_X2 U684 ( .B1(n899), .B2(U1_C_16_), .A(n900), .ZN(n898) );
  AND2_X1 U685 ( .A1(U1_C_15_), .A2(n1464), .ZN(n446) );
  OAI21_X2 U686 ( .B1(n1562), .B2(n65), .A(n980), .ZN(n929) );
  OAI21_X2 U690 ( .B1(U1_C_17_), .B2(n933), .A(U1_C_18_), .ZN(n980) );
  AOI21_X2 U691 ( .B1(n1008), .B2(n609), .A(n1540), .ZN(n958) );
  OAI21_X2 U692 ( .B1(n609), .B2(n1008), .A(U1_C_20_), .ZN(n1039) );
  AOI21_X2 U693 ( .B1(n1038), .B2(n1036), .A(n1543), .ZN(n991) );
  OAI21_X2 U697 ( .B1(n1036), .B2(n1038), .A(n41), .ZN(n1055) );
  AOI21_X2 U700 ( .B1(n1053), .B2(n1051), .A(n1544), .ZN(n1048) );
  OAI21_X2 U701 ( .B1(n1051), .B2(n1053), .A(n29), .ZN(n1088) );
  OAI21_X2 U702 ( .B1(n1554), .B2(n41), .A(n1070), .ZN(n1022) );
  OAI21_X2 U703 ( .B1(U1_C_21_), .B2(n1071), .A(U1_C_22_), .ZN(n1070) );
  OAI21_X2 U704 ( .B1(n1549), .B2(n29), .A(n1099), .ZN(n1080) );
  OAI21_X2 U705 ( .B1(U1_C_23_), .B2(n1084), .A(U1_C_24_), .ZN(n1099) );
  AOI21_X2 U706 ( .B1(n1077), .B2(n1075), .A(n1545), .ZN(n1095) );
  OAI21_X2 U707 ( .B1(n1075), .B2(n1077), .A(n18), .ZN(n1113) );
  OAI21_X2 U708 ( .B1(U1_C_27_), .B2(n368), .A(U1_C_28_), .ZN(n367) );
  OAI21_X2 U709 ( .B1(n1108), .B2(n1110), .A(n12), .ZN(n1122) );
  OAI21_X2 U710 ( .B1(U1_C_25_), .B2(n1093), .A(U1_C_26_), .ZN(n1117) );
  INV_X4 U711 ( .A(n508), .ZN(n208) );
  NAND2_X1 U712 ( .A1(n456), .A2(n277), .ZN(n600) );
  OAI22_X1 U714 ( .A1(n456), .A2(n605), .B1(n619), .B2(n277), .ZN(n606) );
  OAI22_X1 U715 ( .A1(n644), .A2(n277), .B1(n456), .B2(n619), .ZN(n623) );
  OAI22_X1 U716 ( .A1(n456), .A2(n1465), .B1(n474), .B2(n277), .ZN(n471) );
  OAI22_X1 U718 ( .A1(n456), .A2(n644), .B1(n1466), .B2(n277), .ZN(n1231) );
  OAI22_X1 U719 ( .A1(n456), .A2(n1466), .B1(n1465), .B2(n277), .ZN(n1472) );
  OAI22_X1 U720 ( .A1(n456), .A2(n474), .B1(n492), .B2(n277), .ZN(n477) );
  OAI22_X1 U721 ( .A1(n456), .A2(n493), .B1(n494), .B2(n277), .ZN(n482) );
  OAI22_X1 U724 ( .A1(n493), .A2(n277), .B1(n456), .B2(n492), .ZN(n1183) );
  OAI22_X1 U725 ( .A1(n456), .A2(n494), .B1(n695), .B2(n235), .ZN(n496) );
  OAI22_X1 U728 ( .A1(n456), .A2(n695), .B1(n716), .B2(n234), .ZN(n1126) );
  XOR2_X2 U730 ( .A(n387), .B(in_m_mac[4]), .Z(n562) );
  XOR2_X1 U731 ( .A(n694), .B(in_m_mac[4]), .Z(n714) );
  XOR2_X1 U732 ( .A(n1468), .B(in_m_mac[15]), .Z(n642) );
  XOR2_X1 U733 ( .A(n1468), .B(in_m_mac[14]), .Z(n640) );
  XOR2_X1 U734 ( .A(n1468), .B(in_m_mac[13]), .Z(n1469) );
  XOR2_X1 U735 ( .A(n1468), .B(in_m_mac[12]), .Z(n1475) );
  XOR2_X1 U736 ( .A(n1468), .B(in_m_mac[11]), .Z(n1474) );
  XOR2_X1 U737 ( .A(n1468), .B(in_m_mac[10]), .Z(n1164) );
  XOR2_X1 U738 ( .A(n1468), .B(in_m_mac[9]), .Z(n1091) );
  XOR2_X1 U739 ( .A(n1468), .B(in_m_mac[8]), .Z(n1074) );
  XOR2_X1 U741 ( .A(n1468), .B(in_m_mac[7]), .Z(n686) );
  XOR2_X1 U742 ( .A(n1468), .B(in_m_mac[6]), .Z(n684) );
  INV_X8 U743 ( .A(n387), .ZN(n461) );
  XOR2_X1 U744 ( .A(n1413), .B(n346), .Z(n258) );
  XOR2_X1 U745 ( .A(n1425), .B(n1424), .Z(n255) );
  XOR2_X1 U746 ( .A(n1510), .B(n373), .Z(n259) );
  NOR2_X1 U747 ( .A1(n773), .A2(n772), .ZN(n785) );
  INV_X1 U748 ( .A(n1519), .ZN(n1520) );
  INV_X4 U751 ( .A(n787), .ZN(n789) );
  XOR2_X1 U752 ( .A(n788), .B(n791), .Z(n595) );
  OAI22_X1 U753 ( .A1(n744), .A2(n691), .B1(n739), .B2(n690), .ZN(n738) );
  XNOR2_X1 U755 ( .A(n1498), .B(n333), .ZN(n274) );
  NOR2_X1 U757 ( .A1(n439), .A2(n219), .ZN(U5_Z_13) );
  NOR2_X1 U758 ( .A1(n439), .A2(n223), .ZN(U5_Z_8) );
  NOR2_X1 U762 ( .A1(n439), .A2(n242), .ZN(U5_Z_12) );
  NOR2_X1 U763 ( .A1(n439), .A2(n245), .ZN(U5_Z_9) );
  NOR2_X1 U766 ( .A1(n439), .A2(n255), .ZN(U5_Z_3) );
  NOR2_X1 U767 ( .A1(n439), .A2(n244), .ZN(U5_Z_10) );
  NOR2_X1 U769 ( .A1(n439), .A2(n250), .ZN(U5_Z_4) );
  NOR2_X1 U771 ( .A1(n247), .A2(n439), .ZN(U5_Z_7) );
  NOR2_X1 U772 ( .A1(n248), .A2(n439), .ZN(U5_Z_6) );
  NOR2_X1 U773 ( .A1(n249), .A2(n439), .ZN(U5_Z_5) );
  NOR2_X1 U774 ( .A1(n257), .A2(n439), .ZN(U5_Z_1) );
  NOR2_X1 U775 ( .A1(n256), .A2(n439), .ZN(U5_Z_2) );
  NOR2_X1 U778 ( .A1(n819), .A2(n808), .ZN(n820) );
  OAI22_X1 U779 ( .A1(n456), .A2(n714), .B1(n754), .B2(n234), .ZN(n683) );
  OAI22_X1 U780 ( .A1(n456), .A2(n716), .B1(n714), .B2(n235), .ZN(n782) );
  XOR2_X1 U782 ( .A(in_m_mac[2]), .B(n1468), .Z(n559) );
  XOR2_X1 U783 ( .A(n320), .B(n1572), .Z(n617) );
  XNOR2_X1 U786 ( .A(n320), .B(n463), .ZN(n692) );
  XOR2_X1 U787 ( .A(n320), .B(n1573), .Z(n757) );
  XOR2_X1 U788 ( .A(in_m_mac[4]), .B(n1572), .Z(n693) );
  XNOR2_X1 U790 ( .A(in_m_mac[4]), .B(n463), .ZN(n758) );
  XOR2_X1 U792 ( .A(in_m_mac[4]), .B(n1573), .Z(n827) );
  INV_X4 U793 ( .A(n840), .ZN(n448) );
  INV_X1 U798 ( .A(n1491), .ZN(n1493) );
  XNOR2_X1 U799 ( .A(n1415), .B(n293), .ZN(n1417) );
  XOR2_X1 U802 ( .A(n295), .B(n1438), .Z(n1441) );
  INV_X1 U803 ( .A(n1439), .ZN(n1322) );
  XOR2_X1 U804 ( .A(n290), .B(n1434), .Z(n1437) );
  INV_X1 U805 ( .A(n1435), .ZN(n1310) );
  XOR2_X1 U806 ( .A(n291), .B(n1446), .Z(n1449) );
  INV_X1 U807 ( .A(n1447), .ZN(n1349) );
  XNOR2_X1 U808 ( .A(in_m_mac[1]), .B(n463), .ZN(n641) );
  XOR2_X1 U812 ( .A(n356), .B(n1573), .Z(n725) );
  XOR2_X1 U813 ( .A(n356), .B(n1574), .Z(n813) );
  XOR2_X1 U814 ( .A(n356), .B(n1575), .Z(n872) );
  INV_X1 U815 ( .A(n563), .ZN(n449) );
  INV_X1 U816 ( .A(n327), .ZN(n450) );
  INV_X4 U817 ( .A(n450), .ZN(n451) );
  XNOR2_X1 U818 ( .A(n267), .B(n531), .ZN(n522) );
  INV_X4 U820 ( .A(n452), .ZN(n453) );
  XOR2_X1 U821 ( .A(n1457), .B(n265), .Z(n243) );
  INV_X1 U824 ( .A(n1502), .ZN(n454) );
  XOR2_X1 U825 ( .A(n345), .B(n1573), .Z(n822) );
  XOR2_X1 U826 ( .A(n345), .B(n1575), .Z(n943) );
  XOR2_X1 U827 ( .A(n345), .B(n1574), .Z(n875) );
  XNOR2_X1 U828 ( .A(n345), .B(n463), .ZN(n723) );
  XNOR2_X1 U829 ( .A(n284), .B(n261), .ZN(n534) );
  XNOR2_X1 U830 ( .A(n1421), .B(n348), .ZN(n256) );
  XNOR2_X1 U832 ( .A(n1453), .B(n358), .ZN(n244) );
  XNOR2_X1 U833 ( .A(n1429), .B(n453), .ZN(n250) );
  AOI21_X1 U835 ( .B1(n246), .B2(n468), .A(n1090), .ZN(n1086) );
  OAI22_X1 U840 ( .A1(n468), .A2(n1090), .B1(n1063), .B2(n246), .ZN(n1053) );
  OAI22_X1 U841 ( .A1(n468), .A2(n1063), .B1(n1056), .B2(n246), .ZN(n1062) );
  OAI22_X1 U842 ( .A1(n468), .A2(n1056), .B1(n1040), .B2(n246), .ZN(n1036) );
  OAI22_X1 U843 ( .A1(n468), .A2(n1040), .B1(n1012), .B2(n246), .ZN(n1008) );
  OAI22_X1 U848 ( .A1(n468), .A2(n981), .B1(n950), .B2(n246), .ZN(n933) );
  OAI22_X1 U850 ( .A1(n468), .A2(n1012), .B1(n981), .B2(n246), .ZN(n974) );
  OAI22_X1 U851 ( .A1(n468), .A2(n950), .B1(n901), .B2(n246), .ZN(n948) );
  OAI22_X1 U852 ( .A1(n468), .A2(n901), .B1(n874), .B2(n246), .ZN(n855) );
  OAI22_X1 U853 ( .A1(n468), .A2(n874), .B1(n830), .B2(n246), .ZN(n801) );
  OAI22_X1 U854 ( .A1(n468), .A2(n830), .B1(n817), .B2(n246), .ZN(n784) );
  XOR2_X1 U856 ( .A(in_z_mac[7]), .B(in_z_mac[6]), .Z(n1067) );
  INV_X1 U857 ( .A(n636), .ZN(n502) );
  XOR2_X1 U858 ( .A(n1468), .B(in_m_mac[3]), .Z(n582) );
  XOR2_X1 U863 ( .A(n272), .B(n1486), .Z(n1488) );
  NAND2_X1 U864 ( .A1(n590), .A2(n334), .ZN(n594) );
  NAND2_X4 U865 ( .A1(n1067), .A2(n455), .ZN(n1462) );
  INV_X4 U867 ( .A(n470), .ZN(n485) );
  XOR2_X2 U869 ( .A(n694), .B(in_m_mac[11]), .Z(n1465) );
  INV_X4 U870 ( .A(n471), .ZN(n487) );
  NOR2_X2 U875 ( .A1(n471), .A2(n470), .ZN(n473) );
  XOR2_X2 U876 ( .A(n1464), .B(U1_C_15_), .Z(n486) );
  INV_X4 U879 ( .A(n486), .ZN(n472) );
  OAI22_X2 U880 ( .A1(n485), .A2(n487), .B1(n473), .B2(n472), .ZN(n765) );
  INV_X4 U881 ( .A(n477), .ZN(n479) );
  INV_X4 U882 ( .A(n784), .ZN(n475) );
  NOR2_X2 U883 ( .A1(n479), .A2(n475), .ZN(n476) );
  OAI22_X2 U885 ( .A1(n784), .A2(n477), .B1(n476), .B2(n478), .ZN(n824) );
  INV_X4 U887 ( .A(n639), .ZN(n635) );
  INV_X4 U888 ( .A(n1190), .ZN(n701) );
  NOR2_X2 U889 ( .A1(n699), .A2(n701), .ZN(n480) );
  OR2_X1 U890 ( .A1(n777), .A2(n480), .ZN(n736) );
  OAI22_X2 U893 ( .A1(n748), .A2(n322), .B1(n697), .B2(n302), .ZN(n507) );
  NAND2_X2 U894 ( .A1(U1_C_11_), .A2(n507), .ZN(n1144) );
  INV_X4 U899 ( .A(n1144), .ZN(n483) );
  INV_X4 U900 ( .A(n482), .ZN(n1145) );
  NOR2_X2 U901 ( .A1(n1145), .A2(n1144), .ZN(n481) );
  OAI22_X2 U902 ( .A1(n483), .A2(n482), .B1(n481), .B2(n1143), .ZN(n673) );
  OAI22_X2 U903 ( .A1(n685), .A2(n687), .B1(n484), .B2(n1168), .ZN(n674) );
  XOR2_X2 U906 ( .A(n486), .B(n485), .Z(n488) );
  XOR2_X2 U907 ( .A(n488), .B(n487), .Z(n734) );
  OAI22_X2 U908 ( .A1(n818), .A2(n322), .B1(n747), .B2(n302), .ZN(n1480) );
  XOR2_X2 U910 ( .A(n1480), .B(U1_C_13_), .Z(n1184) );
  NAND2_X2 U911 ( .A1(n459), .A2(n444), .ZN(n490) );
  INV_X4 U912 ( .A(n490), .ZN(n506) );
  NOR2_X2 U913 ( .A1(n490), .A2(n489), .ZN(n491) );
  OAI22_X2 U914 ( .A1(n747), .A2(n322), .B1(n748), .B2(n302), .ZN(n505) );
  OAI22_X2 U918 ( .A1(U1_C_12_), .A2(n506), .B1(n491), .B2(n505), .ZN(n1185)
         );
  INV_X4 U922 ( .A(n1183), .ZN(n1188) );
  INV_X4 U925 ( .A(n496), .ZN(n1119) );
  OAI22_X2 U926 ( .A1(n654), .A2(n496), .B1(n495), .B2(n1107), .ZN(n647) );
  OR2_X1 U929 ( .A1(n715), .A2(n497), .ZN(n708) );
  OAI22_X2 U930 ( .A1(n697), .A2(n322), .B1(n661), .B2(n302), .ZN(n501) );
  INV_X4 U931 ( .A(n705), .ZN(n500) );
  INV_X4 U935 ( .A(n501), .ZN(n706) );
  NOR2_X2 U936 ( .A1(n706), .A2(n498), .ZN(n499) );
  OAI22_X2 U938 ( .A1(U1_C_10_), .A2(n501), .B1(n500), .B2(n499), .ZN(n624) );
  NOR2_X2 U942 ( .A1(n713), .A2(n502), .ZN(n503) );
  OAI22_X2 U945 ( .A1(n693), .A2(n455), .B1(n666), .B2(n1462), .ZN(n712) );
  INV_X4 U947 ( .A(n1147), .ZN(n645) );
  OR4_X1 U949 ( .A1(sendz_count[1]), .A2(sendz_count[0]), .A3(n294), .A4(
        sendz_count[2]), .ZN(n508) );
  XOR2_X2 U950 ( .A(n514), .B(U1_C_0_), .Z(n509) );
  NOR2_X2 U951 ( .A1(n208), .A2(n509), .ZN(U6_Z_0) );
  NAND2_X2 U952 ( .A1(n510), .A2(U1_C_1_), .ZN(n520) );
  NOR2_X2 U953 ( .A1(n301), .A2(n458), .ZN(n512) );
  NAND2_X2 U954 ( .A1(n516), .A2(n515), .ZN(n521) );
  NOR3_X2 U955 ( .A1(n517), .A2(n349), .A3(n208), .ZN(U6_Z_1) );
  OAI22_X2 U956 ( .A1(n528), .A2(n322), .B1(n518), .B2(n746), .ZN(n533) );
  NAND2_X2 U957 ( .A1(n521), .A2(n520), .ZN(n531) );
  NOR2_X2 U958 ( .A1(n208), .A2(n522), .ZN(U6_Z_2) );
  NAND2_X2 U959 ( .A1(n386), .A2(n458), .ZN(n523) );
  NAND2_X2 U960 ( .A1(n523), .A2(n364), .ZN(n524) );
  NAND2_X2 U961 ( .A1(n525), .A2(n386), .ZN(n526) );
  XNOR2_X2 U962 ( .A(n537), .B(n541), .ZN(n530) );
  XNOR2_X2 U963 ( .A(n530), .B(n536), .ZN(n548) );
  NOR2_X2 U964 ( .A1(n208), .A2(n535), .ZN(U6_Z_3) );
  INV_X4 U965 ( .A(n536), .ZN(n540) );
  OAI22_X2 U966 ( .A1(n542), .A2(n251), .B1(n540), .B2(n539), .ZN(n569) );
  OAI22_X2 U967 ( .A1(n562), .A2(n322), .B1(n544), .B2(n240), .ZN(n565) );
  NAND2_X2 U968 ( .A1(n546), .A2(n260), .ZN(n547) );
  NOR2_X2 U969 ( .A1(n208), .A2(n550), .ZN(U6_Z_4) );
  NOR2_X2 U970 ( .A1(n336), .A2(n551), .ZN(n552) );
  OAI22_X2 U971 ( .A1(n560), .A2(n322), .B1(n562), .B2(n240), .ZN(n580) );
  OAI22_X2 U972 ( .A1(U1_C_4_), .A2(n449), .B1(n422), .B2(n564), .ZN(n584) );
  INV_X4 U973 ( .A(n569), .ZN(n567) );
  NAND2_X2 U974 ( .A1(n566), .A2(n567), .ZN(n572) );
  NAND2_X2 U975 ( .A1(n568), .A2(n569), .ZN(n570) );
  NAND2_X2 U976 ( .A1(n570), .A2(n218), .ZN(n571) );
  NAND2_X2 U977 ( .A1(n571), .A2(n572), .ZN(n592) );
  NOR2_X2 U978 ( .A1(n208), .A2(n573), .ZN(U6_Z_5) );
  OAI22_X2 U979 ( .A1(n579), .A2(n578), .B1(n576), .B2(n366), .ZN(n828) );
  OAI22_X2 U980 ( .A1(n575), .A2(n322), .B1(n560), .B2(n240), .ZN(n867) );
  NAND2_X2 U981 ( .A1(U1_C_5_), .A2(n580), .ZN(n833) );
  INV_X4 U982 ( .A(n852), .ZN(n835) );
  XNOR2_X2 U983 ( .A(n583), .B(n835), .ZN(n808) );
  INV_X4 U984 ( .A(n584), .ZN(n586) );
  INV_X4 U985 ( .A(n786), .ZN(n791) );
  INV_X4 U986 ( .A(n588), .ZN(n590) );
  NAND2_X2 U987 ( .A1(n594), .A2(n593), .ZN(n787) );
  NOR2_X2 U988 ( .A1(n208), .A2(n598), .ZN(U6_Z_6) );
  INV_X4 U989 ( .A(n1547), .ZN(n1033) );
  XOR2_X2 U990 ( .A(n694), .B(in_m_mac[15]), .Z(n605) );
  INV_X4 U991 ( .A(n605), .ZN(n599) );
  NAND2_X2 U992 ( .A1(n600), .A2(n599), .ZN(n603) );
  INV_X4 U993 ( .A(n603), .ZN(n1279) );
  INV_X4 U994 ( .A(n1004), .ZN(n601) );
  NOR2_X2 U995 ( .A1(n1279), .A2(n601), .ZN(n602) );
  OAI22_X2 U996 ( .A1(n1004), .A2(n603), .B1(n602), .B2(n1278), .ZN(n957) );
  NOR2_X2 U997 ( .A1(n958), .A2(n957), .ZN(n604) );
  OR2_X1 U998 ( .A1(n1035), .A2(n604), .ZN(n994) );
  INV_X4 U999 ( .A(n606), .ZN(n616) );
  INV_X4 U1000 ( .A(n613), .ZN(n608) );
  NOR2_X2 U1001 ( .A1(n52), .A2(n606), .ZN(n607) );
  OAI22_X2 U1002 ( .A1(n616), .A2(n609), .B1(n608), .B2(n607), .ZN(n965) );
  NAND2_X2 U1003 ( .A1(n966), .A2(n965), .ZN(n610) );
  NAND2_X2 U1004 ( .A1(n1013), .A2(n610), .ZN(n1539) );
  INV_X4 U1005 ( .A(n940), .ZN(n612) );
  NOR2_X2 U1006 ( .A1(n940), .A2(n983), .ZN(n611) );
  OAI22_X2 U1007 ( .A1(n612), .A2(n1565), .B1(n1463), .B2(n611), .ZN(n927) );
  XOR2_X2 U1008 ( .A(n613), .B(n609), .Z(n618) );
  XOR2_X2 U1009 ( .A(n618), .B(n616), .Z(n1259) );
  INV_X4 U1010 ( .A(n1259), .ZN(n877) );
  INV_X4 U1011 ( .A(n623), .ZN(n631) );
  INV_X4 U1012 ( .A(n936), .ZN(n620) );
  NOR2_X2 U1013 ( .A1(n631), .A2(n620), .ZN(n621) );
  OAI22_X2 U1014 ( .A1(n936), .A2(n623), .B1(n621), .B2(n630), .ZN(n879) );
  INV_X4 U1015 ( .A(n626), .ZN(n1219) );
  INV_X4 U1016 ( .A(n1218), .ZN(n628) );
  NOR2_X2 U1017 ( .A1(n904), .A2(n626), .ZN(n627) );
  OAI22_X2 U1018 ( .A1(n1567), .A2(n1219), .B1(n628), .B2(n627), .ZN(n849) );
  NAND2_X2 U1019 ( .A1(n766), .A2(n765), .ZN(n629) );
  NAND2_X2 U1020 ( .A1(n850), .A2(n629), .ZN(n1529) );
  XOR2_X2 U1021 ( .A(n630), .B(n936), .Z(n632) );
  XOR2_X2 U1022 ( .A(n632), .B(n631), .Z(n1248) );
  INV_X4 U1023 ( .A(n1248), .ZN(n836) );
  INV_X4 U1024 ( .A(n633), .ZN(n638) );
  NOR2_X2 U1025 ( .A1(n635), .A2(n634), .ZN(n637) );
  OAI22_X2 U1026 ( .A1(U1_C_14_), .A2(n639), .B1(n638), .B2(n637), .ZN(n776)
         );
  INV_X4 U1027 ( .A(n649), .ZN(n1232) );
  NOR2_X2 U1028 ( .A1(n1232), .A2(U1_C_17_), .ZN(n646) );
  XOR2_X2 U1029 ( .A(n694), .B(in_m_mac[12]), .Z(n1466) );
  OAI22_X2 U1030 ( .A1(n65), .A2(n649), .B1(n646), .B2(n1231), .ZN(n889) );
  NAND2_X2 U1031 ( .A1(n930), .A2(n927), .ZN(n650) );
  NAND2_X2 U1032 ( .A1(n979), .A2(n650), .ZN(n1536) );
  NOR2_X2 U1033 ( .A1(n880), .A2(n879), .ZN(n651) );
  OR2_X1 U1034 ( .A1(n968), .A2(n651), .ZN(n925) );
  INV_X4 U1035 ( .A(n655), .ZN(n1380) );
  INV_X4 U1036 ( .A(n368), .ZN(n652) );
  XOR2_X2 U1037 ( .A(n652), .B(n1120), .Z(n1379) );
  INV_X4 U1038 ( .A(n1379), .ZN(n659) );
  NAND2_X2 U1039 ( .A1(n1110), .A2(n1108), .ZN(n653) );
  NOR2_X2 U1040 ( .A1(n1379), .A2(n655), .ZN(n656) );
  OAI22_X2 U1041 ( .A1(n1380), .A2(n659), .B1(n226), .B2(n656), .ZN(n1398) );
  OAI22_X2 U1042 ( .A1(n369), .A2(n361), .B1(n363), .B2(n465), .ZN(n1390) );
  NAND2_X2 U1043 ( .A1(n368), .A2(U1_C_27_), .ZN(n660) );
  NAND2_X2 U1044 ( .A1(n367), .A2(n660), .ZN(n1388) );
  INV_X4 U1045 ( .A(n1388), .ZN(n663) );
  XOR2_X2 U1046 ( .A(n1386), .B(n663), .Z(n664) );
  XOR2_X2 U1047 ( .A(n1390), .B(n664), .Z(n1397) );
  NAND2_X2 U1048 ( .A1(n1081), .A2(n1078), .ZN(n667) );
  NAND2_X2 U1049 ( .A1(n1098), .A2(n667), .ZN(n670) );
  INV_X4 U1050 ( .A(n670), .ZN(n1360) );
  INV_X4 U1051 ( .A(n1093), .ZN(n668) );
  XOR2_X2 U1052 ( .A(n668), .B(n1092), .Z(n1359) );
  INV_X4 U1053 ( .A(n1359), .ZN(n672) );
  INV_X4 U1054 ( .A(n1095), .ZN(n669) );
  XOR2_X2 U1055 ( .A(n669), .B(n1094), .Z(n1358) );
  NOR2_X2 U1056 ( .A1(n1359), .A2(n670), .ZN(n671) );
  OAI22_X2 U1057 ( .A1(n1360), .A2(n672), .B1(n1358), .B2(n671), .ZN(n1371) );
  OAI22_X2 U1058 ( .A1(n615), .A2(n322), .B1(n591), .B2(n240), .ZN(n745) );
  INV_X4 U1059 ( .A(n745), .ZN(n679) );
  NOR2_X2 U1060 ( .A1(n679), .A2(n678), .ZN(n680) );
  OAI22_X2 U1061 ( .A1(U1_C_8_), .A2(n745), .B1(n428), .B2(n680), .ZN(n744) );
  INV_X4 U1062 ( .A(n683), .ZN(n937) );
  NOR2_X2 U1063 ( .A1(n937), .A2(n681), .ZN(n682) );
  OAI22_X2 U1064 ( .A1(n617), .A2(n455), .B1(n596), .B2(n1462), .ZN(n934) );
  OAI22_X2 U1065 ( .A1(n935), .A2(n683), .B1(n682), .B2(n934), .ZN(n691) );
  OAI22_X2 U1066 ( .A1(n457), .A2(n686), .B1(n684), .B2(n362), .ZN(n696) );
  OAI22_X2 U1067 ( .A1(n666), .A2(n455), .B1(n617), .B2(n1462), .ZN(n698) );
  INV_X4 U1068 ( .A(n698), .ZN(n704) );
  INV_X4 U1069 ( .A(n691), .ZN(n742) );
  INV_X4 U1070 ( .A(n744), .ZN(n688) );
  NOR2_X2 U1071 ( .A1(n742), .A2(n688), .ZN(n690) );
  INV_X4 U1072 ( .A(n738), .ZN(n729) );
  OAI22_X2 U1073 ( .A1(n661), .A2(n322), .B1(n615), .B2(n302), .ZN(n718) );
  NAND2_X2 U1074 ( .A1(U1_C_9_), .A2(n718), .ZN(n1128) );
  INV_X4 U1075 ( .A(n696), .ZN(n703) );
  NOR2_X2 U1076 ( .A1(n1569), .A2(n698), .ZN(n700) );
  OAI22_X2 U1077 ( .A1(n662), .A2(n704), .B1(n703), .B2(n700), .ZN(n1127) );
  INV_X4 U1078 ( .A(n1127), .ZN(n1130) );
  INV_X4 U1079 ( .A(n720), .ZN(n783) );
  XOR2_X2 U1080 ( .A(n718), .B(U1_C_9_), .Z(n781) );
  OAI22_X2 U1081 ( .A1(n782), .A2(n720), .B1(n719), .B2(n781), .ZN(n1135) );
  INV_X4 U1082 ( .A(n728), .ZN(n735) );
  NOR2_X2 U1083 ( .A1(n735), .A2(n738), .ZN(n724) );
  OAI22_X2 U1084 ( .A1(n729), .A2(n728), .B1(n737), .B2(n724), .ZN(n1490) );
  INV_X4 U1085 ( .A(n739), .ZN(n743) );
  OAI22_X2 U1086 ( .A1(n591), .A2(n322), .B1(n575), .B2(n240), .ZN(n859) );
  NAND2_X2 U1087 ( .A1(n440), .A2(n458), .ZN(n750) );
  INV_X4 U1088 ( .A(n857), .ZN(n760) );
  OAI22_X2 U1089 ( .A1(n596), .A2(n455), .B1(n597), .B2(n1462), .ZN(n759) );
  NOR2_X2 U1090 ( .A1(n858), .A2(n857), .ZN(n756) );
  OAI22_X2 U1091 ( .A1(n760), .A2(n759), .B1(n756), .B2(n856), .ZN(n764) );
  NAND2_X2 U1092 ( .A1(n762), .A2(n764), .ZN(n916) );
  NAND2_X2 U1093 ( .A1(n918), .A2(n916), .ZN(n769) );
  NAND2_X2 U1094 ( .A1(n769), .A2(n915), .ZN(n1016) );
  INV_X4 U1095 ( .A(n1016), .ZN(n772) );
  OAI22_X2 U1096 ( .A1(n262), .A2(n1016), .B1(n785), .B2(n1006), .ZN(n1044) );
  NAND2_X2 U1097 ( .A1(n789), .A2(n791), .ZN(n805) );
  NAND2_X2 U1098 ( .A1(n793), .A2(n805), .ZN(n1513) );
  OAI22_X2 U1099 ( .A1(n829), .A2(n828), .B1(n825), .B2(n820), .ZN(n1514) );
  NAND2_X2 U1100 ( .A1(n1513), .A2(n1514), .ZN(n832) );
  NOR2_X2 U1101 ( .A1(n835), .A2(n833), .ZN(n851) );
  OAI22_X2 U1102 ( .A1(n457), .A2(n864), .B1(n860), .B2(n362), .ZN(n939) );
  INV_X4 U1103 ( .A(n939), .ZN(n962) );
  OAI22_X2 U1104 ( .A1(U1_C_6_), .A2(n867), .B1(n429), .B2(n866), .ZN(n956) );
  INV_X4 U1105 ( .A(n956), .ZN(n951) );
  INV_X4 U1106 ( .A(n907), .ZN(n895) );
  INV_X4 U1107 ( .A(n1514), .ZN(n876) );
  INV_X4 U1108 ( .A(n905), .ZN(n892) );
  NOR2_X2 U1109 ( .A1(n895), .A2(n892), .ZN(n903) );
  INV_X4 U1110 ( .A(n969), .ZN(n1518) );
  NAND2_X2 U1111 ( .A1(n916), .A2(n915), .ZN(n917) );
  XNOR2_X2 U1112 ( .A(n918), .B(n917), .ZN(n1005) );
  NOR2_X2 U1113 ( .A1(n951), .A2(n939), .ZN(n954) );
  INV_X4 U1114 ( .A(n1003), .ZN(n978) );
  NOR2_X2 U1115 ( .A1(n982), .A2(n978), .ZN(n988) );
  OAI22_X2 U1116 ( .A1(n275), .A2(n1003), .B1(n988), .B2(n986), .ZN(n1522) );
  INV_X4 U1117 ( .A(n1006), .ZN(n1015) );
  AOI21_X4 U1118 ( .B1(n1521), .B2(n1522), .A(n1519), .ZN(n1020) );
  INV_X4 U1119 ( .A(n1044), .ZN(n1489) );
  INV_X4 U1120 ( .A(n1045), .ZN(n1486) );
  NOR2_X2 U1121 ( .A1(n1489), .A2(n1486), .ZN(n1041) );
  INV_X4 U1122 ( .A(n1153), .ZN(n1149) );
  INV_X4 U1123 ( .A(n1126), .ZN(n1131) );
  NOR2_X2 U1124 ( .A1(n1127), .A2(n1126), .ZN(n1129) );
  OAI22_X2 U1125 ( .A1(n1131), .A2(n1130), .B1(n1129), .B2(n1128), .ZN(n1148)
         );
  INV_X4 U1126 ( .A(n1148), .ZN(n1154) );
  INV_X4 U1127 ( .A(n1132), .ZN(n1136) );
  NAND2_X2 U1128 ( .A1(n289), .A2(n1490), .ZN(n1137) );
  OAI22_X2 U1129 ( .A1(n398), .A2(n1142), .B1(n1141), .B2(n1140), .ZN(n1156)
         );
  INV_X4 U1130 ( .A(n1156), .ZN(n1495) );
  XOR2_X2 U1131 ( .A(n1144), .B(n1143), .Z(n1146) );
  XNOR2_X2 U1132 ( .A(n1146), .B(n1145), .ZN(n1172) );
  INV_X4 U1133 ( .A(n1157), .ZN(n1163) );
  INV_X4 U1134 ( .A(n1150), .ZN(n1151) );
  INV_X4 U1135 ( .A(n1162), .ZN(n1158) );
  OAI22_X2 U1136 ( .A1(n333), .A2(n1156), .B1(n1155), .B2(n1496), .ZN(n1176)
         );
  NOR2_X2 U1137 ( .A1(n1158), .A2(n1157), .ZN(n1161) );
  INV_X4 U1138 ( .A(n1159), .ZN(n1160) );
  OAI22_X2 U1139 ( .A1(n1163), .A2(n1162), .B1(n1161), .B2(n1160), .ZN(n1175)
         );
  INV_X4 U1140 ( .A(n1175), .ZN(n1500) );
  NOR2_X2 U1141 ( .A1(n1502), .A2(n1500), .ZN(n1174) );
  XOR2_X2 U1142 ( .A(n1477), .B(n755), .Z(n1165) );
  XNOR2_X2 U1143 ( .A(n1165), .B(n752), .ZN(n1189) );
  INV_X4 U1144 ( .A(n675), .ZN(n1166) );
  XOR2_X2 U1145 ( .A(n1166), .B(n676), .Z(n1179) );
  OR2_X1 U1146 ( .A1(n689), .A2(n1167), .ZN(n1170) );
  INV_X4 U1147 ( .A(n1170), .ZN(n1525) );
  XNOR2_X2 U1148 ( .A(n685), .B(n687), .ZN(n1169) );
  XNOR2_X2 U1150 ( .A(n1169), .B(n1168), .ZN(n1171) );
  INV_X4 U1151 ( .A(n1171), .ZN(n1524) );
  NOR2_X2 U1152 ( .A1(n1171), .A2(n1170), .ZN(n1173) );
  OAI22_X2 U1153 ( .A1(n1525), .A2(n1524), .B1(n1173), .B2(n1172), .ZN(n1177)
         );
  OAI22_X2 U1154 ( .A1(n1181), .A2(n1180), .B1(n1179), .B2(n1178), .ZN(n1193)
         );
  INV_X4 U1155 ( .A(n1193), .ZN(n1503) );
  INV_X4 U1156 ( .A(n1505), .ZN(n1182) );
  NOR2_X2 U1157 ( .A1(n1182), .A2(n1503), .ZN(n1192) );
  INV_X4 U1158 ( .A(n1184), .ZN(n1187) );
  NOR2_X2 U1161 ( .A1(n1184), .A2(n1183), .ZN(n1186) );
  OAI22_X2 U1165 ( .A1(n1188), .A2(n1187), .B1(n1186), .B2(n1185), .ZN(n1204)
         );
  OAI22_X2 U1168 ( .A1(n674), .A2(n673), .B1(n751), .B2(n1189), .ZN(n1206) );
  INV_X4 U1169 ( .A(n1206), .ZN(n1203) );
  INV_X4 U1170 ( .A(n1195), .ZN(n1200) );
  NAND2_X2 U1171 ( .A1(n1526), .A2(n708), .ZN(n1191) );
  NAND2_X2 U1172 ( .A1(n707), .A2(n1191), .ZN(n1199) );
  INV_X4 U1173 ( .A(n1199), .ZN(n1194) );
  OAI22_X2 U1174 ( .A1(n375), .A2(n1193), .B1(n1192), .B2(n1504), .ZN(n1209)
         );
  NOR2_X2 U1175 ( .A1(n1195), .A2(n1194), .ZN(n1198) );
  INV_X4 U1176 ( .A(n1196), .ZN(n1197) );
  OAI22_X2 U1177 ( .A1(n1200), .A2(n1199), .B1(n1198), .B2(n1197), .ZN(n1508)
         );
  INV_X4 U1178 ( .A(n730), .ZN(n1201) );
  XOR2_X2 U1179 ( .A(n1201), .B(n731), .Z(n1211) );
  INV_X4 U1180 ( .A(n1211), .ZN(n1216) );
  INV_X4 U1181 ( .A(n380), .ZN(n1202) );
  NOR2_X2 U1182 ( .A1(n1203), .A2(n1202), .ZN(n1205) );
  OAI22_X2 U1183 ( .A1(n380), .A2(n1206), .B1(n1205), .B2(n1204), .ZN(n1215)
         );
  INV_X4 U1184 ( .A(n1215), .ZN(n1210) );
  INV_X4 U1185 ( .A(n1508), .ZN(n1207) );
  NOR2_X2 U1186 ( .A1(n1509), .A2(n1207), .ZN(n1208) );
  NOR2_X2 U1187 ( .A1(n1211), .A2(n1210), .ZN(n1214) );
  INV_X4 U1188 ( .A(n1212), .ZN(n1213) );
  OAI22_X2 U1189 ( .A1(n1216), .A2(n1215), .B1(n1214), .B2(n1213), .ZN(n1224)
         );
  INV_X4 U1190 ( .A(n1224), .ZN(n1410) );
  INV_X4 U1191 ( .A(n1225), .ZN(n1412) );
  NAND2_X2 U1192 ( .A1(n771), .A2(n1217), .ZN(n1226) );
  XOR2_X2 U1193 ( .A(n1218), .B(n1567), .Z(n1220) );
  XOR2_X2 U1194 ( .A(n1220), .B(n1219), .Z(n763) );
  XOR2_X2 U1195 ( .A(n763), .B(n766), .Z(n1221) );
  XNOR2_X2 U1196 ( .A(n1221), .B(n765), .ZN(n1229) );
  INV_X4 U1197 ( .A(n1229), .ZN(n1227) );
  INV_X4 U1198 ( .A(n1411), .ZN(n1222) );
  OAI22_X2 U1199 ( .A1(n298), .A2(n1224), .B1(n1223), .B2(n1222), .ZN(n1414)
         );
  INV_X4 U1200 ( .A(n1226), .ZN(n1230) );
  NOR2_X2 U1201 ( .A1(n1227), .A2(n1226), .ZN(n1228) );
  OAI22_X2 U1202 ( .A1(n1230), .A2(n1229), .B1(n1228), .B2(n414), .ZN(n1239)
         );
  INV_X4 U1203 ( .A(n1239), .ZN(n1416) );
  NOR2_X2 U1204 ( .A1(n1414), .A2(n1416), .ZN(n1238) );
  XNOR2_X2 U1205 ( .A(n792), .B(n790), .ZN(n1234) );
  XOR2_X2 U1206 ( .A(n1231), .B(n65), .Z(n1233) );
  XOR2_X2 U1207 ( .A(n1233), .B(n1232), .Z(n1538) );
  XNOR2_X2 U1208 ( .A(n1234), .B(n1538), .ZN(n1246) );
  INV_X4 U1209 ( .A(n1246), .ZN(n1240) );
  OR2_X1 U1210 ( .A1(n795), .A2(n1236), .ZN(n1245) );
  INV_X4 U1211 ( .A(n1245), .ZN(n1241) );
  INV_X4 U1212 ( .A(n1415), .ZN(n1237) );
  NOR2_X2 U1213 ( .A1(n1241), .A2(n1240), .ZN(n1244) );
  INV_X4 U1214 ( .A(n1242), .ZN(n1243) );
  OAI22_X2 U1215 ( .A1(n1246), .A2(n1245), .B1(n1244), .B2(n1243), .ZN(n1418)
         );
  INV_X4 U1216 ( .A(n1418), .ZN(n1247) );
  NOR2_X2 U1217 ( .A1(n1420), .A2(n1247), .ZN(n1251) );
  XOR2_X2 U1218 ( .A(n1248), .B(n837), .Z(n1257) );
  XOR2_X2 U1219 ( .A(n1257), .B(n1256), .Z(n1249) );
  INV_X4 U1220 ( .A(n1253), .ZN(n1258) );
  XNOR2_X2 U1221 ( .A(n1249), .B(n1258), .ZN(n1419) );
  INV_X4 U1222 ( .A(n1419), .ZN(n1250) );
  OAI22_X2 U1223 ( .A1(n347), .A2(n1418), .B1(n1251), .B2(n1250), .ZN(n1267)
         );
  INV_X4 U1224 ( .A(n1257), .ZN(n1254) );
  NOR2_X2 U1225 ( .A1(n1254), .A2(n1253), .ZN(n1255) );
  OAI22_X2 U1226 ( .A1(n1258), .A2(n1257), .B1(n1256), .B2(n1255), .ZN(n1266)
         );
  INV_X4 U1227 ( .A(n1266), .ZN(n1422) );
  XOR2_X2 U1228 ( .A(n1259), .B(n880), .Z(n1260) );
  XNOR2_X2 U1229 ( .A(n1260), .B(n879), .ZN(n1268) );
  XOR2_X2 U1230 ( .A(n927), .B(n928), .Z(n1276) );
  XOR2_X2 U1231 ( .A(n1276), .B(n882), .Z(n1270) );
  XOR2_X2 U1232 ( .A(n1268), .B(n1270), .Z(n1263) );
  INV_X4 U1233 ( .A(n1538), .ZN(n1261) );
  OR2_X1 U1234 ( .A1(n885), .A2(n1262), .ZN(n1272) );
  INV_X4 U1235 ( .A(n1272), .ZN(n1269) );
  XNOR2_X2 U1236 ( .A(n1263), .B(n1269), .ZN(n1423) );
  INV_X4 U1237 ( .A(n1423), .ZN(n1264) );
  INV_X4 U1238 ( .A(n1268), .ZN(n1273) );
  NOR2_X2 U1239 ( .A1(n1269), .A2(n1268), .ZN(n1271) );
  INV_X4 U1240 ( .A(n1426), .ZN(n1274) );
  INV_X4 U1241 ( .A(n889), .ZN(n1275) );
  INV_X4 U1242 ( .A(n1276), .ZN(n1277) );
  OAI22_X2 U1243 ( .A1(n884), .A2(n1523), .B1(n926), .B2(n1277), .ZN(n1289) );
  XOR2_X2 U1244 ( .A(n965), .B(n964), .Z(n1461) );
  XOR2_X2 U1245 ( .A(n1278), .B(n1004), .Z(n1280) );
  XOR2_X2 U1246 ( .A(n1280), .B(n1279), .Z(n919) );
  XOR2_X2 U1247 ( .A(n919), .B(n920), .Z(n1286) );
  INV_X4 U1248 ( .A(n1286), .ZN(n1288) );
  XOR2_X2 U1249 ( .A(n221), .B(n1288), .Z(n1281) );
  XOR2_X2 U1250 ( .A(n1289), .B(n1281), .Z(n1427) );
  OAI22_X2 U1251 ( .A1(n452), .A2(n1426), .B1(n1283), .B2(n1282), .ZN(n1290)
         );
  INV_X4 U1252 ( .A(n1289), .ZN(n1285) );
  NOR2_X2 U1253 ( .A1(n1286), .A2(n1285), .ZN(n1287) );
  OAI22_X2 U1254 ( .A1(n1289), .A2(n1288), .B1(n221), .B2(n1287), .ZN(n1298)
         );
  INV_X4 U1255 ( .A(n1298), .ZN(n1432) );
  NOR2_X2 U1256 ( .A1(n1290), .A2(n1432), .ZN(n1297) );
  NAND2_X2 U1257 ( .A1(n1536), .A2(n925), .ZN(n1291) );
  NAND2_X2 U1258 ( .A1(n963), .A2(n1291), .ZN(n1302) );
  INV_X4 U1259 ( .A(n959), .ZN(n1292) );
  XOR2_X2 U1260 ( .A(n958), .B(n955), .Z(n1294) );
  INV_X4 U1261 ( .A(n957), .ZN(n1293) );
  XNOR2_X2 U1262 ( .A(n1294), .B(n1293), .ZN(n1299) );
  INV_X4 U1263 ( .A(n1299), .ZN(n1303) );
  XOR2_X2 U1264 ( .A(n224), .B(n1303), .Z(n1295) );
  XOR2_X2 U1265 ( .A(n1302), .B(n1295), .Z(n1431) );
  INV_X4 U1266 ( .A(n1431), .ZN(n1296) );
  OAI22_X2 U1267 ( .A1(n1430), .A2(n1298), .B1(n1297), .B2(n1296), .ZN(n1435)
         );
  INV_X4 U1268 ( .A(n1302), .ZN(n1300) );
  NOR2_X2 U1269 ( .A1(n1300), .A2(n1299), .ZN(n1301) );
  OAI22_X2 U1270 ( .A1(n1303), .A2(n1302), .B1(n1301), .B2(n224), .ZN(n1436)
         );
  INV_X4 U1271 ( .A(n1436), .ZN(n1304) );
  NOR2_X2 U1272 ( .A1(n1435), .A2(n1304), .ZN(n1309) );
  NAND2_X2 U1273 ( .A1(n1539), .A2(n997), .ZN(n1305) );
  NAND2_X2 U1274 ( .A1(n996), .A2(n1305), .ZN(n1314) );
  INV_X4 U1275 ( .A(n992), .ZN(n1306) );
  INV_X4 U1276 ( .A(n989), .ZN(n1307) );
  XOR2_X2 U1277 ( .A(n1307), .B(n990), .Z(n1315) );
  INV_X4 U1278 ( .A(n1315), .ZN(n1311) );
  XOR2_X2 U1279 ( .A(n225), .B(n1311), .Z(n1308) );
  XOR2_X2 U1280 ( .A(n1314), .B(n1308), .Z(n1434) );
  OAI22_X2 U1281 ( .A1(n1310), .A2(n1436), .B1(n1309), .B2(n1434), .ZN(n1439)
         );
  INV_X4 U1282 ( .A(n1314), .ZN(n1312) );
  NOR2_X2 U1283 ( .A1(n1312), .A2(n1311), .ZN(n1313) );
  OAI22_X2 U1284 ( .A1(n1315), .A2(n1314), .B1(n1313), .B2(n225), .ZN(n1440)
         );
  INV_X4 U1285 ( .A(n1440), .ZN(n1316) );
  INV_X4 U1286 ( .A(n1022), .ZN(n1317) );
  XOR2_X2 U1287 ( .A(n1317), .B(n1021), .Z(n1324) );
  INV_X4 U1288 ( .A(n1025), .ZN(n1318) );
  XOR2_X2 U1289 ( .A(n1318), .B(n1026), .Z(n1326) );
  XOR2_X2 U1290 ( .A(n1324), .B(n1326), .Z(n1320) );
  NAND2_X2 U1291 ( .A1(n995), .A2(n994), .ZN(n1319) );
  NAND2_X2 U1292 ( .A1(n1029), .A2(n1319), .ZN(n1323) );
  INV_X4 U1293 ( .A(n1323), .ZN(n1328) );
  XNOR2_X2 U1294 ( .A(n1320), .B(n1328), .ZN(n1438) );
  OAI22_X2 U1295 ( .A1(n1322), .A2(n1440), .B1(n1321), .B2(n1438), .ZN(n1335)
         );
  INV_X4 U1296 ( .A(n1324), .ZN(n1327) );
  NOR2_X2 U1297 ( .A1(n1324), .A2(n1323), .ZN(n1325) );
  OAI22_X2 U1298 ( .A1(n1328), .A2(n1327), .B1(n1326), .B2(n1325), .ZN(n1443)
         );
  NAND2_X2 U1299 ( .A1(n1028), .A2(n1027), .ZN(n1329) );
  NAND2_X2 U1300 ( .A1(n1050), .A2(n1329), .ZN(n1336) );
  INV_X4 U1301 ( .A(n1046), .ZN(n1330) );
  XOR2_X2 U1302 ( .A(n1330), .B(n1047), .Z(n1338) );
  INV_X4 U1303 ( .A(n1338), .ZN(n1341) );
  NAND2_X2 U1304 ( .A1(n1023), .A2(n1022), .ZN(n1331) );
  NAND2_X2 U1305 ( .A1(n1068), .A2(n1331), .ZN(n1337) );
  INV_X4 U1306 ( .A(n1337), .ZN(n1342) );
  XOR2_X2 U1307 ( .A(n1341), .B(n1342), .Z(n1332) );
  XOR2_X2 U1308 ( .A(n1336), .B(n1332), .Z(n1442) );
  INV_X4 U1309 ( .A(n1443), .ZN(n1333) );
  INV_X4 U1310 ( .A(n1335), .ZN(n1444) );
  OAI22_X2 U1311 ( .A1(n370), .A2(n1443), .B1(n1334), .B2(n1442), .ZN(n1447)
         );
  INV_X4 U1312 ( .A(n1336), .ZN(n1340) );
  NOR2_X2 U1313 ( .A1(n1338), .A2(n1337), .ZN(n1339) );
  OAI22_X2 U1314 ( .A1(n1342), .A2(n1341), .B1(n1340), .B2(n1339), .ZN(n1348)
         );
  INV_X4 U1315 ( .A(n1348), .ZN(n1448) );
  NOR2_X2 U1316 ( .A1(n1447), .A2(n1448), .ZN(n1347) );
  INV_X4 U1317 ( .A(n1078), .ZN(n1343) );
  XOR2_X2 U1318 ( .A(n1343), .B(n1079), .Z(n1352) );
  INV_X4 U1319 ( .A(n1075), .ZN(n1344) );
  XOR2_X2 U1320 ( .A(n1344), .B(n1076), .Z(n1351) );
  INV_X4 U1321 ( .A(n1351), .ZN(n1356) );
  XOR2_X2 U1322 ( .A(n1352), .B(n1356), .Z(n1346) );
  NOR2_X2 U1323 ( .A1(n1049), .A2(n1048), .ZN(n1345) );
  OR2_X1 U1324 ( .A1(n1082), .A2(n1345), .ZN(n1355) );
  INV_X4 U1325 ( .A(n1355), .ZN(n1350) );
  XOR2_X2 U1326 ( .A(n1346), .B(n1350), .Z(n1446) );
  OAI22_X2 U1327 ( .A1(n1349), .A2(n1348), .B1(n1347), .B2(n1446), .ZN(n1363)
         );
  NOR2_X2 U1328 ( .A1(n1351), .A2(n1350), .ZN(n1354) );
  INV_X4 U1329 ( .A(n1352), .ZN(n1353) );
  OAI22_X2 U1330 ( .A1(n1356), .A2(n1355), .B1(n1354), .B2(n1353), .ZN(n1451)
         );
  INV_X4 U1331 ( .A(n1451), .ZN(n1357) );
  INV_X4 U1332 ( .A(n1363), .ZN(n1452) );
  XOR2_X2 U1333 ( .A(n1359), .B(n1358), .Z(n1361) );
  XNOR2_X2 U1334 ( .A(n1361), .B(n1360), .ZN(n1450) );
  INV_X4 U1335 ( .A(n1370), .ZN(n1456) );
  INV_X4 U1336 ( .A(n1371), .ZN(n1454) );
  INV_X4 U1337 ( .A(n1108), .ZN(n1364) );
  XOR2_X2 U1338 ( .A(n1364), .B(n1109), .Z(n1372) );
  INV_X4 U1339 ( .A(n1097), .ZN(n1553) );
  NOR2_X2 U1340 ( .A1(n1095), .A2(n1553), .ZN(n1365) );
  OR2_X1 U1341 ( .A1(n1111), .A2(n1365), .ZN(n1374) );
  XOR2_X2 U1342 ( .A(n1372), .B(n1374), .Z(n1367) );
  NAND2_X2 U1343 ( .A1(n1093), .A2(U1_C_25_), .ZN(n1366) );
  NAND2_X2 U1344 ( .A1(n1117), .A2(n1366), .ZN(n1376) );
  INV_X4 U1345 ( .A(n1376), .ZN(n1373) );
  XNOR2_X2 U1346 ( .A(n1367), .B(n1373), .ZN(n1455) );
  INV_X4 U1347 ( .A(n1455), .ZN(n1368) );
  OAI22_X2 U1348 ( .A1(n1371), .A2(n297), .B1(n1369), .B2(n1368), .ZN(n1384)
         );
  INV_X4 U1349 ( .A(n1372), .ZN(n1377) );
  NOR2_X2 U1350 ( .A1(n1373), .A2(n1372), .ZN(n1375) );
  OAI22_X2 U1351 ( .A1(n1377), .A2(n1376), .B1(n1375), .B2(n1374), .ZN(n1458)
         );
  INV_X4 U1352 ( .A(n1458), .ZN(n1378) );
  XOR2_X2 U1353 ( .A(n1379), .B(n226), .Z(n1381) );
  XOR2_X2 U1354 ( .A(n1381), .B(n1380), .Z(n1459) );
  INV_X4 U1355 ( .A(n1459), .ZN(n1382) );
  NOR2_X2 U1356 ( .A1(n208), .A2(n219), .ZN(U6_Z_29) );
  INV_X4 U1357 ( .A(n1390), .ZN(n1387) );
  NOR2_X2 U1358 ( .A1(n1387), .A2(n1386), .ZN(n1389) );
  OAI22_X2 U1359 ( .A1(n4), .A2(n1390), .B1(n1389), .B2(n1388), .ZN(n1401) );
  NAND2_X2 U1360 ( .A1(n361), .A2(n465), .ZN(n1392) );
  INV_X4 U1361 ( .A(n363), .ZN(n1391) );
  NAND2_X2 U1362 ( .A1(n1392), .A2(n1391), .ZN(n1406) );
  XOR2_X2 U1363 ( .A(U1_C_30_), .B(n1386), .Z(n1393) );
  XOR2_X2 U1364 ( .A(n1406), .B(n1393), .Z(n1400) );
  INV_X4 U1365 ( .A(n1400), .ZN(n1404) );
  INV_X4 U1366 ( .A(n1398), .ZN(n1395) );
  NOR2_X2 U1367 ( .A1(n1394), .A2(n1395), .ZN(n1396) );
  OAI22_X2 U1368 ( .A1(n299), .A2(n1398), .B1(n1396), .B2(n1397), .ZN(n1403)
         );
  NOR2_X2 U1369 ( .A1(n208), .A2(n423), .ZN(U6_Z_30) );
  OAI22_X2 U1370 ( .A1(n1404), .A2(n296), .B1(n1402), .B2(n1401), .ZN(n1409)
         );
  NOR2_X2 U1371 ( .A1(n4), .A2(n1405), .ZN(n1407) );
  OAI22_X2 U1372 ( .A1(U1_C_30_), .A2(n1386), .B1(n1407), .B2(n1406), .ZN(
        n1408) );
  XOR2_X2 U1373 ( .A(n1411), .B(n1410), .Z(n1413) );
  XNOR2_X2 U1374 ( .A(n1417), .B(n1416), .ZN(n257) );
  XNOR2_X2 U1375 ( .A(n1419), .B(n1418), .ZN(n1421) );
  XOR2_X2 U1376 ( .A(n1423), .B(n1422), .Z(n1425) );
  XNOR2_X2 U1377 ( .A(n1427), .B(n1426), .ZN(n1429) );
  XOR2_X2 U1378 ( .A(n1431), .B(n1430), .Z(n1433) );
  XOR2_X2 U1379 ( .A(n1433), .B(n1432), .Z(n249) );
  XNOR2_X2 U1380 ( .A(n1437), .B(n1436), .ZN(n248) );
  XNOR2_X2 U1381 ( .A(n1441), .B(n1440), .ZN(n247) );
  XNOR2_X2 U1382 ( .A(n1449), .B(n1448), .ZN(n245) );
  XOR2_X2 U1383 ( .A(n1451), .B(n1450), .Z(n1453) );
  XOR2_X2 U1384 ( .A(n1455), .B(n1454), .Z(n1457) );
  INV_X4 U1385 ( .A(n1461), .ZN(n923) );
  INV_X4 U1386 ( .A(n1539), .ZN(n961) );
  INV_X4 U1387 ( .A(n997), .ZN(n1541) );
  XOR2_X2 U1388 ( .A(n940), .B(n1463), .Z(n938) );
  INV_X4 U1389 ( .A(n849), .ZN(n1548) );
  OAI22_X2 U1390 ( .A1(n1467), .A2(n1472), .B1(n863), .B2(n865), .ZN(n848) );
  INV_X4 U1391 ( .A(n1481), .ZN(n1471) );
  NOR2_X2 U1392 ( .A1(n1471), .A2(n1470), .ZN(n1552) );
  INV_X4 U1393 ( .A(n1529), .ZN(n846) );
  OAI22_X2 U1394 ( .A1(n1476), .A2(n1482), .B1(n778), .B2(n780), .ZN(n775) );
  INV_X4 U1395 ( .A(n1477), .ZN(n1479) );
  NOR2_X2 U1396 ( .A1(n1479), .A2(n1478), .ZN(n1559) );
  NAND2_X2 U1397 ( .A1(U1_C_13_), .A2(n1480), .ZN(n740) );
  INV_X4 U1398 ( .A(n740), .ZN(n1528) );
  INV_X4 U1399 ( .A(n809), .ZN(n1558) );
  XOR2_X2 U1400 ( .A(n1482), .B(n780), .Z(n779) );
  INV_X4 U1401 ( .A(n1483), .ZN(n1485) );
  NOR2_X2 U1402 ( .A1(n1485), .A2(n1484), .ZN(n1564) );
  XOR2_X2 U1403 ( .A(n1489), .B(n1488), .Z(n283) );
  XNOR2_X2 U1404 ( .A(n1496), .B(n1495), .ZN(n1498) );
  INV_X4 U1405 ( .A(n800), .ZN(n1527) );
  INV_X4 U1406 ( .A(n891), .ZN(n1530) );
  INV_X4 U1407 ( .A(n896), .ZN(n1531) );
  INV_X4 U1408 ( .A(n790), .ZN(n1532) );
  INV_X4 U1409 ( .A(n886), .ZN(n1533) );
  INV_X4 U1410 ( .A(n898), .ZN(n1535) );
  INV_X4 U1411 ( .A(n931), .ZN(n1537) );
  INV_X4 U1412 ( .A(n1039), .ZN(n1540) );
  INV_X4 U1413 ( .A(n1054), .ZN(n1542) );
  INV_X4 U1414 ( .A(n1055), .ZN(n1543) );
  INV_X4 U1415 ( .A(n1088), .ZN(n1544) );
  INV_X4 U1416 ( .A(n1113), .ZN(n1545) );
  INV_X4 U1417 ( .A(n1086), .ZN(n1546) );
  INV_X4 U1418 ( .A(n1084), .ZN(n1549) );
  INV_X4 U1419 ( .A(n1062), .ZN(n1550) );
  INV_X4 U1420 ( .A(n844), .ZN(n1551) );
  INV_X4 U1421 ( .A(n1071), .ZN(n1554) );
  INV_X4 U1422 ( .A(n1058), .ZN(n1555) );
  INV_X4 U1423 ( .A(n1009), .ZN(n1556) );
  INV_X4 U1424 ( .A(n942), .ZN(n1557) );
  INV_X4 U1425 ( .A(n1102), .ZN(n1560) );
  INV_X4 U1426 ( .A(n1032), .ZN(n1561) );
  INV_X4 U1427 ( .A(n933), .ZN(n1562) );
  INV_X4 U1428 ( .A(n948), .ZN(n1563) );
  INV_X4 U1429 ( .A(n983), .ZN(n1565) );
  INV_X4 U1430 ( .A(n871), .ZN(n1566) );
  INV_X4 U1431 ( .A(n904), .ZN(n1567) );
  INV_X4 U1432 ( .A(n812), .ZN(n1568) );
  INV_X4 U1433 ( .A(n662), .ZN(n1569) );
  INV_X4 U1434 ( .A(n710), .ZN(n1570) );
endmodule


module MyDesign ( dut__xxx__finish, xxx__dut__go, dut__bvm__address, 
        dut__bvm__enable, dut__bvm__write, dut__bvm__data, bvm__dut__data, 
        dut__dim__address, dut__dim__enable, dut__dim__write, dut__dim__data, 
        dim__dut__data, dut__dom__address, dut__dom__data, dut__dom__enable, 
        dut__dom__write, clk, reset );
  output [9:0] dut__bvm__address;
  output [15:0] dut__bvm__data;
  input [15:0] bvm__dut__data;
  output [8:0] dut__dim__address;
  output [15:0] dut__dim__data;
  input [15:0] dim__dut__data;
  output [2:0] dut__dom__address;
  output [15:0] dut__dom__data;
  input xxx__dut__go, clk, reset;
  output dut__xxx__finish, dut__bvm__enable, dut__bvm__write, dut__dim__enable,
         dut__dim__write, dut__dom__enable, dut__dom__write;
  wire   n636, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
         n2349, n2350, n2351, n2352, n2353, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
         n2381, n2382, n2383, n2384, n2385, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
         n4888, n4890, n4906, n4910, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n5041, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
         n5056, U8_DATA2_1, U8_DATA2_2, U8_DATA2_3, U8_DATA2_4, U8_DATA2_5,
         U8_DATA2_6, U8_DATA2_7, U8_DATA2_8, U7_DATA2_1, U7_DATA2_2,
         U7_DATA2_3, U7_DATA2_4, U4_DATA1_7, U4_DATA1_8, U4_DATA1_9,
         add_1445_carry_8_, add_1445_B_0_, add_1445_B_1_, add_1445_B_2_,
         add_1445_B_3_, add_1445_B_4_, add_1445_B_5_, add_1445_B_6_,
         add_1445_B_7_, add_1445_B_8_, add_1445_B_9_, add_283_A_0_,
         add_283_A_1_, add_283_A_2_, add_283_A_3_, add_283_A_4_, add_283_A_5_,
         add_180_A_0_, add_180_A_1_, add_180_A_2_, add_180_A_3_, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10092, n10094, n10095, n10096, n10097, n10099,
         n10101, n10102, n10103, n10104, n10106, n10108, n10109, n10110,
         n10111, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10123, n10125, n10126, n10127, n10128, n10130, n10132,
         n10133, n10134, n10135, n10137, n10139, n10140, n10141, n10142,
         n10144, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10158, n10160, n10161, n10162,
         n10163, n10165, n10167, n10168, n10169, n10170, n10172, n10174,
         n10175, n10177, n10178, n10180, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10191, n10193, n10194, n10195,
         n10196, n10198, n10200, n10201, n10202, n10203, n10205, n10207,
         n10208, n10209, n10210, n10212, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10225, n10228, n10231,
         n10233, n10234, n10235, n10236, n10237, n10240, n10243, n10246,
         n10249, n10250, n10251, n10252, n10253, n10254, n10257, n10260,
         n10264, n10267, n10268, n10269, n10270, n10271, n10274, n10277,
         n10280, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10294, n10297, n10300, n10302, n10303, n10304,
         n10305, n10306, n10309, n10312, n10315, n10318, n10319, n10320,
         n10321, n10322, n10323, n10326, n10329, n10333, n10336, n10337,
         n10338, n10339, n10340, n10343, n10346, n10349, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10363,
         n10366, n10369, n10371, n10372, n10373, n10374, n10375, n10378,
         n10381, n10384, n10387, n10388, n10389, n10390, n10391, n10392,
         n10395, n10398, n10402, n10405, n10406, n10407, n10408, n10409,
         n10412, n10415, n10418, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10432, n10435, n10438, n10440,
         n10441, n10442, n10443, n10444, n10447, n10450, n10453, n10456,
         n10457, n10458, n10459, n10460, n10461, n10464, n10467, n10471,
         n10474, n10475, n10476, n10477, n10478, n10481, n10484, n10487,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10501, n10504, n10507, n10509, n10510, n10511, n10512,
         n10513, n10516, n10519, n10522, n10525, n10526, n10527, n10528,
         n10529, n10530, n10533, n10536, n10540, n10543, n10544, n10545,
         n10546, n10547, n10550, n10553, n10556, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10570, n10573,
         n10576, n10578, n10579, n10580, n10581, n10582, n10585, n10588,
         n10591, n10594, n10595, n10596, n10597, n10598, n10599, n10602,
         n10605, n10609, n10612, n10613, n10614, n10615, n10616, n10619,
         n10622, n10625, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10639, n10642, n10645, n10647, n10648,
         n10649, n10650, n10651, n10654, n10657, n10660, n10663, n10664,
         n10665, n10666, n10667, n10668, n10671, n10674, n10678, n10681,
         n10682, n10683, n10684, n10685, n10688, n10691, n10694, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10708, n10711, n10714, n10716, n10717, n10718, n10719, n10720,
         n10723, n10726, n10729, n10732, n10733, n10734, n10735, n10736,
         n10737, n10740, n10743, n10747, n10750, n10751, n10752, n10753,
         n10754, n10757, n10760, n10763, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10777, n10780, n10783,
         n10785, n10786, n10787, n10788, n10789, n10792, n10795, n10798,
         n10801, n10802, n10803, n10804, n10805, n10806, n10809, n10812,
         n10816, n10819, n10820, n10821, n10822, n10823, n10826, n10829,
         n10832, n10836, n10837, n10838, n10839, n10840, n10841, n10842,
         n10843, n10846, n10849, n10852, n10854, n10855, n10856, n10857,
         n10858, n10861, n10864, n10867, n10870, n10871, n10872, n10873,
         n10874, n10875, n10878, n10881, n10885, n10888, n10889, n10890,
         n10891, n10892, n10895, n10898, n10901, n10905, n10906, n10907,
         n10908, n10909, n10910, n10911, n10912, n10915, n10918, n10921,
         n10923, n10924, n10925, n10926, n10927, n10930, n10933, n10936,
         n10939, n10940, n10941, n10942, n10943, n10944, n10947, n10950,
         n10954, n10957, n10958, n10959, n10960, n10961, n10964, n10967,
         n10970, n10974, n10975, n10976, n10977, n10978, n10979, n10980,
         n10981, n10984, n10987, n10990, n10992, n10993, n10994, n10995,
         n10996, n10999, n11002, n11005, n11008, n11009, n11010, n11011,
         n11012, n11013, n11016, n11019, n11023, n11026, n11027, n11028,
         n11029, n11030, n11033, n11036, n11039, n11043, n11044, n11045,
         n11046, n11047, n11048, n11049, n11050, n11053, n11056, n11059,
         n11061, n11062, n11063, n11064, n11065, n11068, n11071, n11074,
         n11077, n11078, n11079, n11080, n11081, n11082, n11085, n11088,
         n11092, n11095, n11096, n11097, n11098, n11099, n11102, n11105,
         n11108, n11112, n11113, n11114, n11115, n11116, n11117, n11118,
         n11119, n11122, n11125, n11128, n11130, n11131, n11132, n11133,
         n11134, n11137, n11140, n11143, n11146, n11147, n11148, n11149,
         n11150, n11151, n11154, n11157, n11161, n11164, n11165, n11166,
         n11167, n11168, n11171, n11174, n11177, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11191, n11192, n11194,
         n11195, n11196, n11199, n11200, n11202, n11203, n11206, n11207,
         n11209, n11212, n11213, n11214, n11215, n11216, n11219, n11220,
         n11221, n11224, n11225, n11226, n11227, n11230, n11231, n11234,
         n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11244,
         n11245, n11246, n11250, n11254, n11257, n11258, n11259, n11260,
         n11261, n11262, n11265, n11266, n11267, n11272, n11275, n11276,
         n11278, n11283, n11399, n11400, n11402, n11419, n11422, n11425,
         n11428, n11430, n11433, n11434, n11435, n11436, n11437, n11438,
         n11439, n11440, n11441, n11452, n11453, n11455, n11457, n11459,
         n11461, n11462, n11464, n11466, n11468, n11470, n11471, n11473,
         n11475, n11477, n11479, n11480, n11482, n11484, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11494, n11496, n11497,
         n11498, n11500, n11501, n11503, n11505, n11507, n11509, n11510,
         n11512, n11514, n11516, n11518, n11519, n11521, n11523, n11525,
         n11527, n11528, n11530, n11532, n11534, n11536, n11537, n11539,
         n11541, n11543, n11545, n11546, n11548, n11550, n11552, n11554,
         n11555, n11557, n11559, n11561, n11563, n11564, n11566, n11568,
         n11570, n11572, n11573, n11575, n11577, n11579, n11581, n11582,
         n11584, n11586, n11588, n11590, n11591, n11593, n11595, n11597,
         n11599, n11600, n11602, n11604, n11606, n11608, n11609, n11611,
         n11613, n11615, n11617, n11618, n11620, n11622, n11624, n11626,
         n11627, n11629, n11631, n11633, n11634, n11636, n11637, n11638,
         n11639, n11640, n11641, n11643, n11645, n11647, n11648, n11649,
         n11651, n11653, n11654, n11655, n11659, n11662, n11663, n11664,
         n11668, n11671, n11672, n11673, n11677, n11680, n11681, n11682,
         n11686, n11689, n11690, n11691, n11695, n11698, n11699, n11700,
         n11704, n11707, n11708, n11709, n11713, n11716, n11717, n11718,
         n11722, n11725, n11726, n11727, n11731, n11734, n11735, n11736,
         n11740, n11743, n11744, n11745, n11749, n11752, n11753, n11754,
         n11758, n11761, n11762, n11763, n11767, n11770, n11771, n11772,
         n11776, n11779, n11780, n11781, n11788, n11789, n11793, n11794,
         n11798, n11801, n11803, n11806, n11809, n11811, n11813, n11815,
         n11874, n11876, n11878, n11880, n12056, n12057, n12058, n12060,
         n12062, n12140, n12145, n12146, n12152, n12153, n12154, n12155,
         n12156, n12157, n12158, n12159, n12160, n12162, n12164, n12165,
         n12167, n12169, n12170, n12172, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12182, n12183, n12185, n12186, n12187,
         n12188, n12190, n12192, n12193, n12194, n12195, n12196, n12197,
         n12198, n12199, n12200, n12201, n12203, n12205, n12207, n12208,
         n12210, n12212, n12213, n12214, n12215, n12216, n12218, n12219,
         n12221, n12223, n12224, n12226, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12237, n12242, n12243, n12246, n12249,
         n12250, n12251, n12252, n12253, n12257, n12260, n12264, n12267,
         n12268, n12269, n12270, n12271, n12272, n12273, n12276, n12281,
         n12282, n12285, n12288, n12289, n12290, n12291, n12292, n12296,
         n12299, n12303, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12315, n12320, n12321, n12324, n12327, n12328, n12329,
         n12330, n12331, n12335, n12338, n12342, n12346, n12347, n12348,
         n12349, n12350, n12351, n12354, n12359, n12360, n12363, n12366,
         n12367, n12368, n12369, n12370, n12374, n12377, n12381, n12385,
         n12386, n12387, n12388, n12389, n12390, n12393, n12398, n12399,
         n12402, n12405, n12406, n12407, n12408, n12409, n12413, n12416,
         n12420, n12424, n12425, n12426, n12427, n12428, n12429, n12432,
         n12437, n12438, n12441, n12444, n12445, n12446, n12447, n12448,
         n12452, n12455, n12459, n12463, n12464, n12465, n12466, n12467,
         n12468, n12471, n12476, n12477, n12480, n12483, n12484, n12485,
         n12486, n12487, n12491, n12494, n12498, n12502, n12503, n12504,
         n12505, n12506, n12507, n12510, n12515, n12516, n12519, n12522,
         n12523, n12524, n12525, n12526, n12530, n12533, n12537, n12541,
         n12542, n12543, n12544, n12545, n12546, n12549, n12554, n12555,
         n12558, n12561, n12562, n12563, n12564, n12565, n12569, n12572,
         n12576, n12580, n12581, n12582, n12583, n12584, n12585, n12588,
         n12593, n12594, n12597, n12600, n12601, n12602, n12603, n12604,
         n12608, n12611, n12615, n12619, n12620, n12621, n12622, n12623,
         n12624, n12627, n12632, n12633, n12636, n12639, n12640, n12641,
         n12642, n12643, n12647, n12650, n12654, n12658, n12659, n12660,
         n12661, n12662, n12663, n12666, n12671, n12672, n12675, n12678,
         n12679, n12680, n12681, n12682, n12686, n12689, n12693, n12697,
         n12698, n12699, n12700, n12701, n12702, n12705, n12710, n12711,
         n12714, n12717, n12718, n12719, n12720, n12721, n12725, n12728,
         n12732, n12736, n12737, n12738, n12739, n12740, n12741, n12744,
         n12749, n12750, n12753, n12756, n12757, n12758, n12759, n12760,
         n12764, n12767, n12771, n12775, n12776, n12777, n12778, n12779,
         n12780, n12783, n12786, n12787, n12788, n12789, n12790, n12791,
         n12794, n12796, n12799, n12800, n12803, n12804, n12805, n12806,
         n12807, n12808, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12820, n12823, n12825, n12826, n12827, n12828, n12829,
         n12830, n12831, n12832, n12835, n12838, n12839, n12840, n12841,
         n12843, n12844, n12846, n12847, n12849, n12853, n12872, n12889,
         n12892, n12910, n12927, n12930, n12948, n12965, n12966, n12967,
         n12968, n12969, n12970, n12971, n12972, n12974, n12975, n12977,
         n12978, n12980, n12982, n12984, n12986, n12988, n12992, n13009,
         n13012, n13029, n13031, n13032, n13043, n13045, n13046, n13050,
         n13051, n13052, n13053, n13054, n13055, n13057, n13058, n13059,
         n13060, n13063, n13065, n13066, n13067, n13068, n13069, n13071,
         n13072, n13073, n13075, n13076, n13077, n13078, n13080, n13081,
         n13083, n13084, n13085, n13086, n13088, n13091, n13092, n13093,
         n13095, n13096, n13099, n13100, n13101, n13102, n13103, n13104,
         n13109, n13119, n13124, n13132, n13137, n13138, n13139, n13140,
         n13144, n13155, n13160, n13166, n13172, n13173, n13174, n13175,
         n13176, n13177, n13180, n13185, n13186, n13189, n13192, n13193,
         n13194, n13195, n13197, n13203, n13204, n13205, n13209, n13210,
         n13211, n13212, n13213, n13214, n13217, n13222, n13223, n13226,
         n13229, n13230, n13231, n13232, n13234, n13240, n13241, n13242,
         n13246, n13247, n13248, n13249, n13250, n13251, n13254, n13259,
         n13260, n13263, n13266, n13267, n13268, n13269, n13271, n13277,
         n13278, n13279, n13283, n13284, n13285, n13286, n13287, n13288,
         n13291, n13296, n13297, n13300, n13303, n13304, n13305, n13306,
         n13308, n13314, n13315, n13316, n13320, n13321, n13322, n13323,
         n13324, n13325, n13328, n13333, n13334, n13337, n13340, n13341,
         n13342, n13343, n13345, n13351, n13352, n13353, n13357, n13358,
         n13359, n13360, n13361, n13362, n13365, n13370, n13371, n13374,
         n13377, n13378, n13379, n13380, n13382, n13388, n13389, n13390,
         n13394, n13395, n13396, n13397, n13398, n13399, n13402, n13407,
         n13408, n13411, n13414, n13415, n13416, n13417, n13419, n13425,
         n13426, n13427, n13431, n13432, n13433, n13434, n13435, n13436,
         n13439, n13444, n13445, n13448, n13451, n13452, n13453, n13454,
         n13456, n13462, n13463, n13464, n13468, n13469, n13470, n13471,
         n13472, n13473, n13476, n13481, n13482, n13485, n13488, n13489,
         n13490, n13491, n13493, n13499, n13500, n13501, n13505, n13506,
         n13507, n13508, n13509, n13510, n13513, n13518, n13519, n13522,
         n13525, n13526, n13527, n13528, n13530, n13536, n13537, n13538,
         n13542, n13543, n13544, n13545, n13546, n13547, n13550, n13555,
         n13556, n13559, n13562, n13563, n13564, n13565, n13567, n13573,
         n13574, n13575, n13578, n13579, n13580, n13581, n13582, n13583,
         n13584, n13587, n13592, n13593, n13596, n13599, n13600, n13601,
         n13602, n13604, n13610, n13611, n13612, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13624, n13629, n13630, n13633,
         n13636, n13637, n13638, n13639, n13641, n13647, n13648, n13649,
         n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13661,
         n13666, n13667, n13670, n13673, n13674, n13675, n13676, n13678,
         n13684, n13685, n13686, n13689, n13690, n13691, n13692, n13693,
         n13694, n13695, n13698, n13703, n13704, n13707, n13710, n13711,
         n13712, n13713, n13715, n13721, n13722, n13723, n13727, n13728,
         n13729, n13730, n13731, n13732, n13735, n13740, n13741, n13744,
         n13747, n13748, n13749, n13750, n13752, n13758, n13759, n13760,
         n13764, n13765, n13766, n13767, n13768, n13769, n13772, n13777,
         n13778, n13781, n13784, n13785, n13786, n13787, n13789, n13795,
         n13796, n13797, n13801, n13802, n13803, n13804, n13805, n13806,
         n13809, n13814, n13815, n13818, n13821, n13822, n13823, n13824,
         n13826, n13832, n13833, n13834, n13838, n13839, n13840, n13841,
         n13842, n13843, n13846, n13851, n13852, n13855, n13858, n13859,
         n13860, n13861, n13863, n13869, n13870, n13871, n13875, n13876,
         n13877, n13878, n13879, n13880, n13883, n13888, n13889, n13892,
         n13895, n13896, n13897, n13898, n13900, n13906, n13907, n13908,
         n13912, n13913, n13914, n13915, n13916, n13917, n13920, n13925,
         n13926, n13929, n13932, n13933, n13934, n13935, n13937, n13943,
         n13944, n13945, n13949, n13950, n13951, n13952, n13953, n13954,
         n13957, n13962, n13963, n13966, n13969, n13970, n13971, n13972,
         n13974, n13980, n13981, n13982, n13986, n13987, n13988, n13989,
         n13990, n13991, n13994, n13999, n14000, n14003, n14006, n14007,
         n14008, n14009, n14011, n14017, n14018, n14019, n14023, n14024,
         n14025, n14026, n14027, n14028, n14031, n14036, n14037, n14040,
         n14043, n14044, n14045, n14046, n14048, n14054, n14055, n14056,
         n14060, n14061, n14062, n14063, n14064, n14065, n14068, n14073,
         n14074, n14077, n14080, n14081, n14082, n14083, n14085, n14091,
         n14092, n14093, n14097, n14098, n14099, n14100, n14101, n14102,
         n14105, n14110, n14111, n14114, n14117, n14118, n14119, n14120,
         n14122, n14128, n14129, n14130, n14134, n14135, n14136, n14137,
         n14138, n14139, n14142, n14147, n14148, n14151, n14154, n14155,
         n14156, n14157, n14159, n14165, n14166, n14167, n14170, n14171,
         n14172, n14173, n14174, n14175, n14176, n14179, n14184, n14185,
         n14188, n14191, n14192, n14193, n14194, n14196, n14202, n14203,
         n14204, n14207, n14208, n14209, n14210, n14211, n14212, n14213,
         n14216, n14221, n14222, n14225, n14228, n14229, n14230, n14231,
         n14233, n14239, n14240, n14241, n14244, n14245, n14246, n14247,
         n14248, n14249, n14250, n14253, n14258, n14259, n14262, n14265,
         n14266, n14267, n14268, n14270, n14276, n14277, n14278, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14290, n14295,
         n14296, n14299, n14302, n14303, n14304, n14305, n14307, n14313,
         n14314, n14315, n14319, n14320, n14321, n14322, n14323, n14324,
         n14327, n14332, n14333, n14336, n14339, n14340, n14341, n14342,
         n14344, n14350, n14351, n14352, n14356, n14357, n14358, n14359,
         n14360, n14361, n14364, n14369, n14370, n14373, n14376, n14377,
         n14378, n14379, n14381, n14387, n14388, n14389, n14393, n14394,
         n14395, n14396, n14397, n14398, n14401, n14406, n14407, n14410,
         n14413, n14414, n14415, n14416, n14418, n14424, n14425, n14426,
         n14430, n14431, n14432, n14433, n14434, n14435, n14438, n14443,
         n14444, n14447, n14450, n14451, n14452, n14453, n14455, n14461,
         n14462, n14463, n14467, n14468, n14469, n14470, n14471, n14472,
         n14475, n14480, n14481, n14484, n14487, n14488, n14489, n14490,
         n14492, n14498, n14499, n14500, n14504, n14505, n14506, n14507,
         n14508, n14509, n14512, n14517, n14518, n14521, n14524, n14525,
         n14526, n14527, n14529, n14535, n14536, n14537, n14541, n14542,
         n14543, n14544, n14545, n14546, n14549, n14554, n14555, n14558,
         n14561, n14562, n14563, n14564, n14566, n14572, n14573, n14574,
         n14578, n14579, n14580, n14581, n14582, n14583, n14586, n14591,
         n14592, n14595, n14598, n14599, n14600, n14601, n14603, n14609,
         n14610, n14611, n14615, n14616, n14617, n14618, n14619, n14620,
         n14623, n14628, n14629, n14632, n14635, n14636, n14637, n14638,
         n14640, n14646, n14647, n14648, n14652, n14653, n14654, n14655,
         n14656, n14657, n14660, n14665, n14666, n14669, n14672, n14673,
         n14674, n14675, n14677, n14683, n14684, n14685, n14689, n14690,
         n14691, n14692, n14693, n14694, n14697, n14702, n14703, n14706,
         n14709, n14710, n14711, n14712, n14714, n14720, n14721, n14722,
         n14726, n14727, n14728, n14729, n14730, n14731, n14734, n14739,
         n14740, n14743, n14746, n14747, n14748, n14749, n14751, n14757,
         n14758, n14759, n14762, n14763, n14764, n14765, n14766, n14767,
         n14768, n14771, n14776, n14777, n14780, n14783, n14784, n14785,
         n14786, n14788, n14794, n14795, n14796, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14808, n14813, n14814, n14817,
         n14820, n14821, n14822, n14823, n14825, n14831, n14832, n14833,
         n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14845,
         n14850, n14851, n14854, n14857, n14858, n14859, n14860, n14862,
         n14868, n14869, n14870, n14873, n14874, n14875, n14876, n14877,
         n14878, n14879, n14882, n14887, n14888, n14891, n14894, n14895,
         n14896, n14897, n14899, n14905, n14906, n14907, n14911, n14912,
         n14913, n14914, n14915, n14916, n14919, n14924, n14925, n14928,
         n14931, n14932, n14933, n14934, n14936, n14942, n14943, n14944,
         n14948, n14949, n14950, n14951, n14952, n14953, n14956, n14961,
         n14962, n14965, n14968, n14969, n14970, n14971, n14973, n14979,
         n14980, n14981, n14985, n14986, n14987, n14988, n14989, n14990,
         n14993, n14998, n14999, n15002, n15005, n15006, n15007, n15008,
         n15010, n15016, n15017, n15018, n15022, n15023, n15024, n15025,
         n15026, n15027, n15030, n15035, n15036, n15039, n15042, n15043,
         n15044, n15045, n15047, n15053, n15054, n15055, n15059, n15060,
         n15061, n15062, n15063, n15064, n15067, n15072, n15073, n15076,
         n15079, n15080, n15081, n15082, n15084, n15090, n15091, n15092,
         n15096, n15097, n15098, n15099, n15100, n15101, n15104, n15109,
         n15110, n15113, n15116, n15117, n15118, n15119, n15121, n15127,
         n15128, n15129, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15141, n15146, n15147, n15150, n15153, n15154, n15155,
         n15156, n15158, n15164, n15165, n15166, n15169, n15170, n15171,
         n15172, n15173, n15174, n15175, n15178, n15183, n15184, n15187,
         n15190, n15191, n15192, n15193, n15195, n15201, n15202, n15203,
         n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15215,
         n15220, n15221, n15224, n15227, n15228, n15229, n15230, n15232,
         n15238, n15239, n15240, n15243, n15244, n15245, n15246, n15247,
         n15248, n15249, n15252, n15257, n15258, n15261, n15264, n15265,
         n15266, n15267, n15269, n15275, n15276, n15277, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15289, n15294, n15295,
         n15298, n15301, n15302, n15303, n15304, n15306, n15312, n15313,
         n15314, n15317, n15318, n15319, n15320, n15321, n15322, n15323,
         n15326, n15331, n15332, n15335, n15338, n15339, n15340, n15341,
         n15343, n15349, n15350, n15351, n15354, n15355, n15356, n15357,
         n15358, n15359, n15360, n15363, n15368, n15369, n15372, n15375,
         n15376, n15377, n15378, n15380, n15386, n15387, n15388, n15391,
         n15392, n15393, n15394, n15395, n15396, n15397, n15400, n15405,
         n15406, n15409, n15412, n15413, n15414, n15415, n15417, n15423,
         n15424, n15425, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15437, n15442, n15443, n15446, n15449, n15450, n15451,
         n15452, n15454, n15460, n15461, n15462, n15465, n15466, n15467,
         n15468, n15469, n15470, n15471, n15474, n15477, n15478, n15479,
         n15480, n15483, n15484, n15485, n15488, n15489, n15492, n15493,
         n15494, n15495, n15497, n15503, n15504, n15505, n15509, n15511,
         n15513, n15514, n15515, n15516, n15517, n15518, n15521, n15522,
         n15523, n15526, n15530, n15531, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15543, n15545, n15546, n15550,
         n15567, n15569, n15572, n15590, n15606, n15609, n15626, n15628,
         n15631, n15649, n15667, n15684, n15686, n15689, n15707, n15741,
         n15743, n15746, n15764, n15780, n15782, n15785, n15803, n15820,
         n15822, n15823, n15825, n15828, n15846, n15863, n15865, n15867,
         n15870, n15888, n15905, n15907, n15909, n15912, n15930, n15947,
         n15949, n15950, n15952, n15955, n15972, n15974, n15976, n15977,
         n15979, n15982, n15999, n16001, n16003, n16005, n16008, n16025,
         n16027, n16029, n16031, n16034, n16051, n16053, n16055, n16059,
         n16076, n16078, n16081, n16099, n16115, n16118, n16135, n16137,
         n16140, n16158, n16174, n16175, n16176, n16177, n16178, n16179,
         n16180, n16181, n16182, n16185, n16188, n16189, n16191, n16192,
         n16193, n16194, n16196, n16199, n16200, n16201, n16202, n16205,
         n16207, n16208, n16209, n16210, n16211, n16216, n16218, n16221,
         n16238, n16240, n16243, n16261, n16279, n16296, n16298, n16300,
         n16303, n16321, n16339, n16341, n16342, n16343, n16344, n16346,
         n16347, n16348, n16351, n16352, n16353, n16354, n16358, n16359,
         n16360, n16361, n16364, n16365, n16366, n16367, n16368, n16369,
         n16370, n16371, n16372, n16373, n16374, n16377, n16378, n16379,
         n16381, n16382, n16383, n16386, n16387, n16390, n16391, n16392,
         n16393, n16394, n16395, n16396, n16398, n16400, n16401, n16402,
         n16403, n16404, n16405, n16407, n16409, n16410, n16411, n16414,
         n16415, n16416, n16418, n16419, n16420, n16423, n16424, n16427,
         n16428, n16429, n16430, n16431, n16432, n16433, n16435, n16437,
         n16438, n16439, n16440, n16441, n16442, n16444, n16446, n16447,
         n16448, n16451, n16452, n16453, n16455, n16456, n16457, n16460,
         n16461, n16464, n16465, n16466, n16467, n16468, n16469, n16470,
         n16472, n16474, n16475, n16476, n16477, n16478, n16479, n16481,
         n16483, n16484, n16485, n16488, n16489, n16490, n16492, n16493,
         n16494, n16497, n16498, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16509, n16511, n16512, n16513, n16514, n16515,
         n16516, n16518, n16520, n16521, n16522, n16525, n16526, n16527,
         n16529, n16530, n16531, n16534, n16535, n16538, n16539, n16540,
         n16541, n16542, n16543, n16544, n16546, n16548, n16549, n16550,
         n16551, n16552, n16553, n16555, n16557, n16558, n16559, n16562,
         n16563, n16564, n16566, n16567, n16568, n16571, n16572, n16575,
         n16576, n16577, n16578, n16579, n16580, n16581, n16583, n16585,
         n16586, n16587, n16588, n16589, n16590, n16592, n16594, n16595,
         n16596, n16599, n16600, n16601, n16603, n16604, n16605, n16608,
         n16609, n16612, n16613, n16614, n16615, n16616, n16617, n16618,
         n16620, n16622, n16623, n16624, n16625, n16626, n16627, n16629,
         n16631, n16632, n16633, n16636, n16637, n16638, n16640, n16641,
         n16642, n16645, n16646, n16649, n16650, n16651, n16652, n16653,
         n16654, n16655, n16657, n16659, n16660, n16661, n16662, n16663,
         n16664, n16666, n16668, n16669, n16670, n16673, n16674, n16675,
         n16677, n16678, n16679, n16682, n16683, n16686, n16687, n16688,
         n16689, n16690, n16691, n16692, n16694, n16696, n16697, n16698,
         n16699, n16700, n16701, n16703, n16705, n16706, n16707, n16710,
         n16711, n16712, n16714, n16715, n16716, n16719, n16720, n16723,
         n16724, n16725, n16726, n16727, n16728, n16729, n16731, n16733,
         n16734, n16735, n16736, n16737, n16738, n16740, n16742, n16743,
         n16744, n16747, n16748, n16749, n16751, n16752, n16753, n16756,
         n16757, n16760, n16761, n16762, n16763, n16764, n16765, n16766,
         n16768, n16770, n16771, n16772, n16773, n16774, n16775, n16777,
         n16779, n16780, n16781, n16784, n16785, n16786, n16788, n16789,
         n16790, n16793, n16794, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16805, n16807, n16808, n16809, n16810, n16811,
         n16812, n16814, n16816, n16817, n16818, n16821, n16822, n16823,
         n16825, n16826, n16827, n16830, n16831, n16834, n16835, n16836,
         n16837, n16838, n16839, n16840, n16842, n16844, n16845, n16846,
         n16847, n16848, n16849, n16851, n16853, n16854, n16855, n16858,
         n16859, n16860, n16862, n16863, n16864, n16867, n16868, n16871,
         n16872, n16873, n16874, n16875, n16876, n16877, n16879, n16881,
         n16882, n16883, n16884, n16885, n16886, n16888, n16890, n16891,
         n16892, n16895, n16896, n16897, n16899, n16900, n16901, n16904,
         n16905, n16908, n16909, n16910, n16911, n16912, n16913, n16914,
         n16916, n16918, n16919, n16920, n16921, n16922, n16923, n16925,
         n16927, n16928, n16929, n16932, n16933, n16934, n16936, n16937,
         n16938, n16941, n16942, n16945, n16946, n16947, n16948, n16949,
         n16950, n16951, n16953, n16955, n16956, n16957, n16958, n16959,
         n16960, n16962, n16964, n16965, n16966, n16969, n16970, n16971,
         n16973, n16974, n16975, n16978, n16979, n16982, n16983, n16984,
         n16985, n16986, n16987, n16988, n16990, n16992, n16993, n16994,
         n16995, n16996, n16997, n16999, n17001, n17002, n17003, n17006,
         n17007, n17008, n17010, n17011, n17012, n17015, n17016, n17019,
         n17020, n17021, n17022, n17023, n17024, n17025, n17027, n17029,
         n17030, n17031, n17032, n17033, n17034, n17036, n17038, n17039,
         n17040, n17043, n17044, n17045, n17047, n17048, n17049, n17052,
         n17053, n17056, n17057, n17058, n17059, n17060, n17061, n17062,
         n17064, n17066, n17067, n17068, n17069, n17070, n17071, n17073,
         n17075, n17076, n17077, n17080, n17081, n17082, n17084, n17085,
         n17086, n17089, n17090, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17101, n17103, n17104, n17105, n17106, n17107,
         n17108, n17110, n17112, n17113, n17114, n17117, n17118, n17119,
         n17121, n17122, n17123, n17126, n17127, n17130, n17131, n17132,
         n17133, n17134, n17135, n17136, n17138, n17140, n17141, n17142,
         n17143, n17144, n17145, n17147, n17149, n17150, n17151, n17154,
         n17155, n17156, n17158, n17159, n17160, n17163, n17164, n17167,
         n17168, n17169, n17170, n17171, n17172, n17173, n17175, n17177,
         n17178, n17179, n17180, n17181, n17182, n17184, n17186, n17187,
         n17188, n17191, n17192, n17193, n17195, n17196, n17197, n17200,
         n17201, n17204, n17205, n17206, n17207, n17208, n17209, n17210,
         n17212, n17214, n17215, n17216, n17217, n17218, n17219, n17221,
         n17223, n17224, n17225, n17228, n17229, n17230, n17232, n17233,
         n17234, n17237, n17238, n17241, n17242, n17243, n17244, n17245,
         n17246, n17247, n17249, n17251, n17252, n17253, n17254, n17255,
         n17256, n17258, n17260, n17261, n17262, n17265, n17266, n17267,
         n17269, n17270, n17271, n17274, n17275, n17278, n17279, n17280,
         n17281, n17282, n17283, n17284, n17286, n17288, n17289, n17290,
         n17291, n17292, n17293, n17295, n17297, n17298, n17299, n17302,
         n17303, n17304, n17306, n17307, n17308, n17311, n17312, n17315,
         n17316, n17317, n17318, n17319, n17320, n17321, n17323, n17325,
         n17326, n17327, n17328, n17329, n17330, n17332, n17334, n17335,
         n17336, n17339, n17340, n17341, n17343, n17344, n17345, n17348,
         n17349, n17352, n17353, n17354, n17355, n17356, n17357, n17358,
         n17360, n17362, n17363, n17364, n17365, n17366, n17367, n17369,
         n17371, n17372, n17373, n17376, n17377, n17378, n17380, n17381,
         n17382, n17385, n17386, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17397, n17399, n17400, n17401, n17402, n17403,
         n17404, n17406, n17408, n17409, n17410, n17413, n17414, n17415,
         n17417, n17418, n17419, n17422, n17423, n17426, n17427, n17428,
         n17429, n17430, n17431, n17432, n17434, n17436, n17437, n17438,
         n17439, n17440, n17441, n17443, n17445, n17446, n17447, n17450,
         n17451, n17452, n17454, n17455, n17456, n17459, n17460, n17463,
         n17464, n17465, n17466, n17467, n17468, n17469, n17471, n17473,
         n17474, n17475, n17476, n17477, n17478, n17480, n17482, n17483,
         n17484, n17487, n17488, n17489, n17491, n17492, n17493, n17496,
         n17497, n17500, n17501, n17502, n17503, n17504, n17505, n17506,
         n17508, n17510, n17511, n17512, n17513, n17514, n17515, n17517,
         n17519, n17520, n17521, n17524, n17525, n17526, n17528, n17529,
         n17530, n17533, n17534, n17537, n17538, n17539, n17540, n17541,
         n17542, n17543, n17545, n17547, n17548, n17549, n17550, n17551,
         n17552, n17554, n17556, n17557, n17558, n17561, n17562, n17563,
         n17565, n17566, n17567, n17570, n17571, n17574, n17575, n17576,
         n17577, n17578, n17579, n17580, n17582, n17584, n17585, n17586,
         n17587, n17588, n17589, n17591, n17593, n17594, n17595, n17598,
         n17599, n17600, n17602, n17603, n17604, n17607, n17608, n17611,
         n17612, n17613, n17614, n17615, n17616, n17617, n17619, n17621,
         n17622, n17623, n17624, n17625, n17626, n17628, n17630, n17631,
         n17632, n17635, n17636, n17637, n17639, n17640, n17641, n17644,
         n17645, n17648, n17649, n17650, n17651, n17652, n17653, n17654,
         n17656, n17658, n17659, n17660, n17661, n17662, n17663, n17665,
         n17667, n17668, n17669, n17672, n17673, n17674, n17676, n17677,
         n17678, n17681, n17682, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17693, n17695, n17696, n17697, n17698, n17699,
         n17700, n17702, n17704, n17705, n17706, n17709, n17710, n17711,
         n17713, n17714, n17715, n17718, n17719, n17722, n17723, n17724,
         n17725, n17726, n17727, n17728, n17730, n17732, n17733, n17734,
         n17735, n17736, n17737, n17739, n17741, n17742, n17743, n17746,
         n17747, n17748, n17750, n17751, n17752, n17755, n17756, n17759,
         n17760, n17761, n17762, n17763, n17764, n17765, n17767, n17769,
         n17770, n17771, n17772, n17773, n17774, n17776, n17778, n17779,
         n17780, n17783, n17784, n17785, n17787, n17788, n17789, n17792,
         n17793, n17796, n17797, n17798, n17799, n17800, n17801, n17802,
         n17804, n17806, n17807, n17808, n17809, n17810, n17811, n17813,
         n17815, n17816, n17817, n17820, n17821, n17822, n17824, n17825,
         n17826, n17829, n17830, n17833, n17834, n17835, n17836, n17837,
         n17838, n17839, n17841, n17843, n17844, n17845, n17846, n17847,
         n17848, n17850, n17852, n17853, n17854, n17857, n17858, n17859,
         n17861, n17862, n17863, n17866, n17867, n17870, n17871, n17872,
         n17873, n17874, n17875, n17876, n17878, n17880, n17881, n17882,
         n17883, n17884, n17885, n17887, n17889, n17890, n17891, n17894,
         n17895, n17896, n17898, n17899, n17900, n17903, n17904, n17907,
         n17908, n17909, n17910, n17911, n17912, n17913, n17915, n17917,
         n17918, n17919, n17920, n17921, n17922, n17924, n17926, n17927,
         n17928, n17931, n17932, n17933, n17935, n17936, n17937, n17940,
         n17941, n17944, n17945, n17946, n17947, n17948, n17949, n17950,
         n17952, n17954, n17955, n17956, n17957, n17958, n17959, n17961,
         n17963, n17964, n17965, n17968, n17969, n17970, n17972, n17973,
         n17974, n17977, n17978, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17989, n17991, n17992, n17993, n17994, n17995,
         n17996, n17998, n18000, n18001, n18002, n18005, n18006, n18007,
         n18009, n18010, n18011, n18014, n18015, n18018, n18019, n18020,
         n18021, n18022, n18023, n18024, n18026, n18028, n18029, n18030,
         n18031, n18032, n18033, n18035, n18037, n18038, n18039, n18042,
         n18043, n18044, n18046, n18047, n18048, n18051, n18052, n18055,
         n18056, n18057, n18058, n18059, n18060, n18061, n18063, n18065,
         n18066, n18067, n18068, n18069, n18070, n18072, n18074, n18075,
         n18076, n18079, n18080, n18081, n18083, n18084, n18085, n18088,
         n18089, n18092, n18093, n18094, n18095, n18096, n18097, n18098,
         n18100, n18102, n18103, n18104, n18105, n18106, n18107, n18109,
         n18111, n18112, n18113, n18116, n18117, n18118, n18120, n18121,
         n18122, n18125, n18126, n18129, n18130, n18131, n18132, n18133,
         n18134, n18135, n18137, n18139, n18140, n18141, n18142, n18143,
         n18144, n18146, n18148, n18149, n18150, n18153, n18154, n18155,
         n18157, n18158, n18159, n18162, n18163, n18166, n18167, n18168,
         n18169, n18170, n18171, n18172, n18174, n18176, n18177, n18178,
         n18179, n18180, n18181, n18183, n18185, n18186, n18187, n18190,
         n18191, n18192, n18194, n18195, n18196, n18199, n18200, n18203,
         n18204, n18205, n18206, n18207, n18208, n18209, n18211, n18213,
         n18214, n18215, n18216, n18217, n18218, n18220, n18222, n18223,
         n18224, n18227, n18228, n18229, n18231, n18232, n18233, n18236,
         n18237, n18240, n18241, n18242, n18243, n18244, n18245, n18246,
         n18248, n18250, n18251, n18252, n18253, n18254, n18255, n18257,
         n18259, n18260, n18261, n18264, n18265, n18266, n18268, n18269,
         n18270, n18273, n18274, n18277, n18278, n18279, n18280, n18281,
         n18282, n18283, n18285, n18287, n18288, n18289, n18290, n18291,
         n18292, n18294, n18296, n18297, n18298, n18301, n18302, n18303,
         n18305, n18306, n18307, n18310, n18311, n18314, n18315, n18316,
         n18317, n18318, n18319, n18320, n18322, n18324, n18325, n18326,
         n18327, n18328, n18329, n18331, n18333, n18334, n18335, n18338,
         n18339, n18340, n18342, n18343, n18344, n18347, n18348, n18351,
         n18352, n18353, n18354, n18355, n18356, n18357, n18359, n18361,
         n18362, n18363, n18364, n18365, n18366, n18368, n18370, n18371,
         n18372, n18375, n18376, n18377, n18379, n18380, n18381, n18384,
         n18385, n18388, n18389, n18390, n18391, n18392, n18393, n18394,
         n18396, n18398, n18399, n18400, n18401, n18402, n18403, n18405,
         n18407, n18408, n18409, n18412, n18413, n18414, n18416, n18417,
         n18418, n18421, n18422, n18425, n18426, n18427, n18428, n18429,
         n18430, n18431, n18433, n18435, n18436, n18437, n18438, n18439,
         n18440, n18442, n18444, n18445, n18446, n18449, n18450, n18451,
         n18453, n18454, n18455, n18458, n18459, n18462, n18463, n18464,
         n18465, n18466, n18467, n18468, n18470, n18472, n18473, n18474,
         n18475, n18476, n18477, n18479, n18481, n18482, n18483, n18486,
         n18487, n18488, n18490, n18491, n18492, n18495, n18496, n18499,
         n18500, n18501, n18502, n18503, n18504, n18505, n18507, n18509,
         n18510, n18511, n18512, n18513, n18514, n18516, n18518, n18519,
         n18520, n18523, n18524, n18525, n18527, n18528, n18529, n18532,
         n18533, n18536, n18537, n18538, n18539, n18540, n18541, n18542,
         n18544, n18546, n18547, n18548, n18549, n18550, n18551, n18553,
         n18555, n18556, n18557, n18560, n18561, n18562, n18564, n18565,
         n18566, n18569, n18570, n18573, n18574, n18575, n18576, n18577,
         n18578, n18579, n18581, n18583, n18584, n18585, n18586, n18587,
         n18588, n18590, n18592, n18593, n18594, n18597, n18598, n18599,
         n18601, n18602, n18603, n18606, n18607, n18610, n18611, n18612,
         n18613, n18614, n18615, n18616, n18618, n18620, n18621, n18622,
         n18623, n18624, n18625, n18627, n18629, n18630, n18631, n18634,
         n18635, n18636, n18638, n18639, n18640, n18643, n18644, n18647,
         n18648, n18649, n18650, n18651, n18652, n18653, n18655, n18657,
         n18658, n18659, n18660, n18661, n18662, n18664, n18666, n18667,
         n18668, n18671, n18672, n18673, n18675, n18676, n18677, n18680,
         n18681, n18684, n18685, n18686, n18687, n18688, n18689, n18690,
         n18692, n18694, n18695, n18696, n18697, n18698, n18699, n18701,
         n18703, n18704, n18705, n18708, n18709, n18710, n18712, n18713,
         n18714, n18717, n18718, n18721, n18722, n18723, n18724, n18725,
         n18726, n18727, n18729, n18731, n18732, n18733, n18734, n18735,
         n18736, n18738, n18740, n18741, n18742, n18743, n18744, n18745,
         n18746, n18747, n18748, n18750, n18751, n18752, n18753, n18754,
         n18755, n18756, n18757, n18758, n18759, n18763, n18764, n18765,
         n18766, n18767, n18768, n18770, n18771, n18772, n18773, n18776,
         n18777, n18781, n18782, n18785, n18786, n18787, n18788, n18790,
         n18791, n18792, n18793, n18794, n18795, n18796, n18800, n18801,
         n18802, n18803, n18804, n18805, n18807, n18808, n18809, n18810,
         n18813, n18814, n18818, n18819, n18822, n18823, n18824, n18825,
         n18827, n18828, n18830, n18831, n18832, n18833, n18837, n18838,
         n18839, n18840, n18841, n18842, n18844, n18845, n18846, n18847,
         n18850, n18851, n18855, n18856, n18859, n18860, n18861, n18862,
         n18864, n18865, n18866, n18867, n18868, n18869, n18870, n18874,
         n18875, n18876, n18877, n18878, n18879, n18881, n18882, n18883,
         n18884, n18887, n18888, n18892, n18893, n18896, n18897, n18898,
         n18899, n18901, n18902, n18903, n18904, n18905, n18906, n18907,
         n18911, n18912, n18913, n18914, n18915, n18916, n18918, n18919,
         n18920, n18921, n18924, n18925, n18929, n18930, n18933, n18934,
         n18935, n18936, n18938, n18939, n18940, n18941, n18942, n18943,
         n18944, n18948, n18949, n18950, n18951, n18952, n18953, n18955,
         n18956, n18957, n18958, n18961, n18962, n18966, n18967, n18970,
         n18971, n18972, n18973, n18975, n18976, n18977, n18978, n18979,
         n18980, n18981, n18985, n18986, n18987, n18988, n18989, n18990,
         n18992, n18993, n18994, n18995, n18998, n18999, n19003, n19004,
         n19007, n19008, n19009, n19010, n19012, n19013, n19014, n19015,
         n19016, n19017, n19018, n19022, n19023, n19024, n19025, n19026,
         n19027, n19029, n19030, n19031, n19032, n19035, n19036, n19040,
         n19041, n19044, n19045, n19046, n19047, n19049, n19050, n19052,
         n19053, n19054, n19055, n19059, n19060, n19061, n19062, n19063,
         n19064, n19066, n19067, n19068, n19069, n19072, n19073, n19077,
         n19078, n19081, n19082, n19083, n19084, n19086, n19087, n19088,
         n19089, n19090, n19091, n19092, n19096, n19097, n19098, n19099,
         n19100, n19101, n19103, n19104, n19105, n19106, n19109, n19110,
         n19114, n19115, n19118, n19119, n19120, n19121, n19123, n19124,
         n19126, n19127, n19128, n19129, n19133, n19134, n19135, n19136,
         n19137, n19138, n19140, n19141, n19142, n19143, n19146, n19147,
         n19151, n19152, n19155, n19156, n19157, n19158, n19160, n19161,
         n19163, n19164, n19165, n19166, n19170, n19171, n19172, n19173,
         n19174, n19175, n19177, n19178, n19179, n19180, n19183, n19184,
         n19188, n19189, n19192, n19193, n19194, n19195, n19197, n19198,
         n19200, n19201, n19202, n19203, n19207, n19208, n19209, n19210,
         n19211, n19212, n19214, n19215, n19216, n19217, n19220, n19221,
         n19225, n19226, n19229, n19230, n19231, n19232, n19234, n19235,
         n19237, n19238, n19239, n19240, n19244, n19245, n19246, n19247,
         n19248, n19249, n19251, n19252, n19253, n19254, n19257, n19258,
         n19262, n19263, n19266, n19267, n19268, n19269, n19271, n19272,
         n19274, n19275, n19276, n19277, n19281, n19282, n19283, n19284,
         n19285, n19286, n19288, n19289, n19290, n19291, n19294, n19295,
         n19299, n19300, n19303, n19304, n19305, n19306, n19308, n19309,
         n19311, n19312, n19313, n19314, n19318, n19319, n19320, n19321,
         n19322, n19323, n19325, n19326, n19327, n19328, n19331, n19332,
         n19336, n19337, n19340, n19341, n19342, n19343, n19345, n19346,
         n19348, n19349, n19350, n19351, n19352, n19355, n19356, n19360,
         n19363, n19364, n19368, n19371, n19372, n19376, n19379, n19380,
         n19384, n19387, n19388, n19392, n19395, n19396, n19400, n19403,
         n19404, n19408, n19411, n19412, n19416, n19419, n19420, n19424,
         n19427, n19428, n19432, n19435, n19436, n19440, n19443, n19444,
         n19448, n19451, n19452, n19456, n19459, n19460, n19464, n19467,
         n19468, n19472, n19475, n19476, n19480, n19481, n19482, n19483,
         n19486, n19487, n19490, n19491, n19492, n19495, n19496, n19499,
         n19500, n19503, n19504, n19507, n19508, n19513, n19514, n19516,
         n19517, n19522, n19523, n19524, n19525, n19530, n19531, n19532,
         n19533, n19538, n19539, n19540, n19541, n19544, n19545, n19547,
         n19548, n19551, n19552, n19555, n19556, n19557, n19560, n19561,
         n19564, n19565, n19568, n19569, n19572, n19573, n19578, n19579,
         n19580, n19581, n19582, n19583, n19584, n19585, n19586, n19587,
         n19588, n19589, n19590, n19591, n19592, n19593, n19594, n19595,
         n19596, n19597, n19598, n19599, n19600, n19601, n19602, n19603,
         n19604, n19605, n19606, n19607, n19608, n19609, n19610, n19611,
         n19612, n19613, n19616, n19617, n19620, n19621, n19622, n19625,
         n19626, n19629, n19630, n19633, n19634, n19637, n19638, n19643,
         n19644, n19645, n19646, n19647, n19648, n19649, n19650, n19651,
         n19652, n19653, n19654, n19655, n19656, n19657, n19658, n19659,
         n19660, n19661, n19662, n19663, n19664, n19665, n19666, n19667,
         n19668, n19669, n19670, n19671, n19672, n19673, n19674, n19675,
         n19676, n19677, n19678, n19681, n19682, n19685, n19686, n19687,
         n19690, n19691, n19694, n19695, n19698, n19699, n19702, n19703,
         n19708, n19709, n19710, n19711, n19712, n19713, n19714, n19715,
         n19716, n19717, n19718, n19719, n19720, n19721, n19722, n19723,
         n19724, n19725, n19726, n19727, n19728, n19729, n19730, n19731,
         n19732, n19733, n19734, n19735, n19736, n19737, n19738, n19739,
         n19740, n19741, n19742, n19743, n19746, n19747, n19750, n19751,
         n19752, n19755, n19756, n19759, n19760, n19763, n19764, n19767,
         n19768, n19773, n19774, n19775, n19776, n19777, n19778, n19779,
         n19780, n19781, n19782, n19783, n19784, n19785, n19786, n19787,
         n19788, n19789, n19790, n19791, n19792, n19793, n19794, n19795,
         n19796, n19797, n19798, n19799, n19800, n19801, n19802, n19803,
         n19804, n19805, n19806, n19807, n19808, n19811, n19812, n19815,
         n19816, n19817, n19820, n19821, n19824, n19825, n19828, n19829,
         n19832, n19833, n19838, n19839, n19840, n19841, n19842, n19843,
         n19844, n19845, n19846, n19847, n19848, n19849, n19850, n19851,
         n19852, n19853, n19854, n19855, n19856, n19857, n19858, n19859,
         n19860, n19861, n19862, n19863, n19864, n19865, n19866, n19867,
         n19868, n19869, n19870, n19871, n19872, n19873, n19876, n19877,
         n19880, n19881, n19882, n19885, n19886, n19889, n19890, n19893,
         n19894, n19897, n19898, n19903, n19904, n19905, n19906, n19907,
         n19908, n19909, n19910, n19911, n19912, n19913, n19914, n19915,
         n19916, n19917, n19918, n19919, n19920, n19921, n19922, n19923,
         n19924, n19925, n19926, n19927, n19928, n19929, n19930, n19931,
         n19932, n19933, n19934, n19935, n19936, n19937, n19938, n19941,
         n19942, n19945, n19946, n19947, n19950, n19951, n19954, n19955,
         n19958, n19959, n19962, n19963, n19968, n19969, n19970, n19971,
         n19972, n19973, n19974, n19975, n19976, n19977, n19978, n19979,
         n19980, n19981, n19982, n19983, n19984, n19985, n19986, n19987,
         n19988, n19989, n19990, n19991, n19992, n19993, n19994, n19995,
         n19996, n19997, n19998, n19999, n20000, n20001, n20002, n20003,
         n20006, n20007, n20010, n20011, n20012, n20015, n20016, n20019,
         n20020, n20023, n20024, n20027, n20028, n20033, n20034, n20035,
         n20036, n20037, n20038, n20039, n20040, n20041, n20042, n20043,
         n20044, n20045, n20046, n20047, n20048, n20049, n20050, n20051,
         n20052, n20053, n20054, n20055, n20056, n20057, n20058, n20059,
         n20060, n20061, n20062, n20063, n20064, n20065, n20066, n20067,
         n20068, n20071, n20072, n20075, n20076, n20077, n20080, n20081,
         n20084, n20085, n20088, n20089, n20092, n20093, n20098, n20099,
         n20100, n20101, n20102, n20103, n20104, n20105, n20106, n20107,
         n20108, n20109, n20110, n20111, n20112, n20113, n20114, n20115,
         n20116, n20117, n20118, n20119, n20120, n20121, n20122, n20123,
         n20124, n20125, n20126, n20127, n20128, n20129, n20130, n20131,
         n20132, n20133, n20136, n20137, n20140, n20141, n20142, n20145,
         n20146, n20149, n20150, n20153, n20154, n20157, n20158, n20163,
         n20164, n20165, n20166, n20167, n20168, n20169, n20170, n20171,
         n20172, n20173, n20174, n20175, n20176, n20177, n20178, n20179,
         n20180, n20181, n20182, n20183, n20184, n20185, n20186, n20187,
         n20188, n20189, n20190, n20191, n20192, n20193, n20194, n20195,
         n20196, n20197, n20198, n20201, n20202, n20205, n20206, n20207,
         n20210, n20211, n20214, n20215, n20218, n20219, n20222, n20223,
         n20228, n20229, n20230, n20231, n20232, n20233, n20234, n20235,
         n20236, n20237, n20238, n20239, n20240, n20241, n20242, n20243,
         n20244, n20245, n20246, n20247, n20248, n20249, n20250, n20251,
         n20252, n20253, n20254, n20255, n20256, n20257, n20258, n20259,
         n20260, n20261, n20262, n20263, n20266, n20267, n20270, n20271,
         n20272, n20275, n20276, n20279, n20280, n20283, n20284, n20287,
         n20288, n20293, n20294, n20295, n20296, n20297, n20298, n20299,
         n20300, n20301, n20302, n20303, n20304, n20305, n20306, n20307,
         n20308, n20309, n20310, n20311, n20312, n20313, n20314, n20315,
         n20316, n20317, n20318, n20319, n20320, n20321, n20322, n20323,
         n20324, n20325, n20326, n20327, n20328, n20331, n20332, n20335,
         n20336, n20337, n20340, n20341, n20344, n20345, n20348, n20349,
         n20352, n20353, n20358, n20359, n20360, n20361, n20362, n20363,
         n20364, n20365, n20366, n20367, n20368, n20369, n20370, n20371,
         n20372, n20373, n20374, n20375, n20376, n20377, n20378, n20379,
         n20380, n20381, n20382, n20383, n20384, n20385, n20386, n20387,
         n20388, n20389, n20390, n20391, n20392, n20393, n20396, n20397,
         n20400, n20401, n20402, n20405, n20406, n20409, n20410, n20413,
         n20414, n20417, n20418, n20423, n20424, n20425, n20426, n20427,
         n20428, n20429, n20430, n20431, n20432, n20433, n20434, n20435,
         n20436, n20437, n20438, n20439, n20440, n20441, n20442, n20443,
         n20444, n20445, n20446, n20447, n20448, n20449, n20450, n20451,
         n20452, n20453, n20454, n20455, n20456, n20457, n20458, n20459,
         n20462, n20463, n20466, n20467, n20468, n20471, n20472, n20475,
         n20476, n20479, n20480, n20483, n20484, n20489, n20490, n20491,
         n20492, n20493, n20494, n20495, n20496, n20497, n20498, n20499,
         n20500, n20501, n20502, n20503, n20504, n20505, n20506, n20507,
         n20508, n20509, n20510, n20511, n20512, n20513, n20514, n20515,
         n20516, n20517, n20518, n20519, n20520, n20521, n20522, n20523,
         n20524, n20525, n20526, n20528, n20529, n20530, n20531, n20532,
         n20533, n20534, n20535, n20536, n20537, n20538, n20539, n20540,
         n20541, n20542, n20543, n20544, n20545, n20546, n20547, n20548,
         n20549, n20550, n20551, n20552, n20553, n20554, n20555, n20556,
         n20557, n20558, n20559, n20560, n20561, n20562, n20563, n20564,
         n20565, n20566, n20567, n20568, n20569, n20570, n20571, n20572,
         n20573, n20574, n20575, n20576, n20577, n20578, n20579, n20580,
         n20581, n20582, n20583, n20584, n20585, n20586, n20588, n20589,
         n20590, n20591, n20592, n20593, n20594, n20595, n20596, n20597,
         n20598, n20599, n20600, n20601, n20602, n20604, n20605, n20606,
         n20607, n20608, n20609, n20610, n20611, n20612, n20613, n20614,
         n20615, n20616, n20617, n20618, n20620, n20621, n20622, n20623,
         n20624, n20625, n20626, n20627, n20628, n20629, n20630, n20631,
         n20632, n20633, n20634, n20636, n20637, n20638, n20639, n20640,
         n20641, n20642, n20643, n20644, n20645, n20646, n20647, n20648,
         n20649, n20650, n20652, n20653, n20654, n20655, n20656, n20657,
         n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665,
         n20666, n20668, n20669, n20670, n20671, n20672, n20673, n20674,
         n20675, n20676, n20677, n20678, n20679, n20680, n20681, n20682,
         n20684, n20685, n20686, n20687, n20688, n20689, n20690, n20691,
         n20692, n20693, n20694, n20695, n20696, n20697, n20698, n20700,
         n20701, n20702, n20703, n20704, n20705, n20706, n20707, n20708,
         n20709, n20710, n20711, n20712, n20713, n20714, n20716, n20717,
         n20718, n20719, n20720, n20721, n20722, n20723, n20724, n20725,
         n20726, n20727, n20728, n20729, n20730, n20732, n20733, n20734,
         n20735, n20736, n20737, n20738, n20739, n20740, n20741, n20742,
         n20743, n20744, n20745, n20746, n20748, n20749, n20750, n20751,
         n20752, n20753, n20754, n20755, n20756, n20757, n20758, n20759,
         n20760, n20761, n20762, n20764, n20765, n20766, n20767, n20768,
         n20769, n20770, n20771, n20772, n20773, n20774, n20775, n20776,
         n20777, n20778, n20780, n20781, n20782, n20783, n20784, n20785,
         n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793,
         n20794, n20796, n20797, n20798, n20799, n20800, n20801, n20802,
         n20803, n20804, n20805, n20806, n20807, n20808, n20809, n20810,
         n20812, n20813, n20814, n20815, n20816, n20817, n20818, n20819,
         n20820, n20821, n20822, n20823, n20824, n20825, n20826, n20828,
         n20829, n20830, n20831, n20832, n20833, n20834, n20835, n20836,
         n20837, n20838, n20839, n20840, n20841, n20842, n20844, n20845,
         n20846, n20847, n20848, n20849, n20850, n20851, n20852, n20853,
         n20854, n20855, n20856, n20857, n20858, n20860, n20861, n20862,
         n20863, n20864, n20865, n20866, n20867, n20868, n20869, n20870,
         n20871, n20872, n20873, n20874, n20876, n20877, n20878, n20879,
         n20880, n20881, n20882, n20883, n20884, n20885, n20886, n20887,
         n20888, n20889, n20890, n20892, n20893, n20894, n20895, n20896,
         n20897, n20898, n20899, n20900, n20901, n20902, n20903, n20904,
         n20905, n20906, n20908, n20909, n20910, n20911, n20912, n20913,
         n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921,
         n20922, n20924, n20925, n20926, n20927, n20928, n20929, n20930,
         n20931, n20932, n20933, n20934, n20935, n20936, n20937, n20938,
         n20940, n20941, n20942, n20943, n20944, n20945, n20946, n20947,
         n20948, n20949, n20950, n20951, n20952, n20953, n20954, n20956,
         n20957, n20958, n20959, n20960, n20961, n20962, n20963, n20964,
         n20965, n20966, n20967, n20968, n20969, n20970, n20972, n20973,
         n20974, n20975, n20976, n20977, n20978, n20979, n20980, n20981,
         n20982, n20983, n20984, n20985, n20986, n20988, n20989, n20990,
         n20991, n20992, n20993, n20994, n20995, n20996, n20997, n20998,
         n20999, n21000, n21001, n21002, n21004, n21005, n21006, n21007,
         n21008, n21009, n21010, n21011, n21012, n21013, n21014, n21015,
         n21016, n21017, n21018, n21020, n21021, n21022, n21023, n21024,
         n21025, n21026, n21027, n21028, n21029, n21030, n21031, n21032,
         n21033, n21034, n21036, n21037, n21038, n21039, n21040, n21041,
         n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049,
         n21050, n21052, n21053, n21054, n21055, n21056, n21057, n21058,
         n21059, n21060, n21061, n21062, n21063, n21064, n21065, n21066,
         n21068, n21069, n21070, n21071, n21072, n21073, n21074, n21075,
         n21076, n21077, n21078, n21079, n21080, n21081, n21082, n21084,
         n21085, n21086, n21087, n21088, n21089, n21090, n21091, n21092,
         n21093, n21094, n21095, n21096, n21097, n21098, n21099, n21100,
         n21101, n21102, n21103, n21104, n21105, n21106, n21107, n21108,
         n21109, n21110, n21111, n21112, n21113, n21114, n21115, n21116,
         n21117, n21118, n21119, n21120, n21121, n21122, n21123, n21124,
         n21125, n21126, n21127, n21128, n21129, n21130, n21131, n21132,
         n21133, n21134, n21135, n21136, n21137, n21138, n21139, n21140,
         n21141, n21142, n21143, n21144, n21145, n21146, n21147, n21148,
         n21149, n21150, n21151, n21152, n21153, n21154, n21155, n21156,
         n21157, n21158, n21159, n21160, n21161, n21162, n21163, n21164,
         n21165, n21166, n21167, n21168, n21169, n21170, n21171, n21172,
         n21173, n21174, n21175, n21176, n21177, n21178, n21179, n21180,
         n21181, n21182, n21183, n21184, n21185, n21186, n21187, n21188,
         n21189, n21190, n21191, n21192, n21193, n21194, n21195, n21196,
         n21197, n21198, n21199, n21200, n21201, n21202, n21203, n21204,
         n21205, n21206, n21207, n21208, n21209, n21210, n21211, n21212,
         n21213, n21214, n21215, n21216, n21217, n21218, n21219, n21220,
         n21221, n21222, n21223, n21224, n21225, n21226, n21227, n21228,
         n21229, n21230, n21231, n21232, n21233, n21234, n21235, n21236,
         n21237, n21238, n21239, n21240, n21241, n21242, n21243, n21244,
         n21245, n21246, n21247, n21248, n21249, n21250, n21251, n21252,
         n21253, n21254, n21255, n21256, n21257, n21258, n21259, n21260,
         n21261, n21262, n21263, n21264, n21265, n21266, n21267, n21268,
         n21269, n21270, n21271, n21272, n21273, n21274, n21275, n21276,
         n21277, n21278, n21279, n21280, n21281, n21282, n21283, n21284,
         n21285, n21286, n21287, n21288, n21289, n21290, n21291, n21292,
         n21293, n21294, n21295, n21296, n21297, n21298, n21299, n21300,
         n21301, n21302, n21303, n21304, n21305, n21306, n21307, n21308,
         n21309, n21310, n21311, n21312, n21313, n21314, n21315, n21316,
         n21317, n21318, n21319, n21320, n21321, n21322, n21323, n21324,
         n21325, n21326, n21327, n21328, n21329, n21330, n21331, n21332,
         n21333, n21334, n21335, n21336, n21337, n21338, n21339, n21340,
         n21341, n21342, n21343, n21344, n21345, n21346, n21347, n21348,
         n21349, n21350, n21351, n21352, n21353, n21354, n21355, n21356,
         n21357, n21358, n21359, n21360, n21361, n21362, n21363, n21364,
         n21365, n21366, n21367, n21368, n21369, n21370, n21371, n21372,
         n21373, n21374, n21375, n21376, n21377, n21378, n21379, n21380,
         n21381, n21382, n21383, n21384, n21385, n21386, n21387, n21388,
         n21389, n21390, n21391, n21392, n21393, n21394, n21395, n21396,
         n21397, n21398, n21399, n21400, n21401, n21402, n21403, n21404,
         n21405, n21406, n21407, n21408, n21409, n21410, n21411, n21412,
         n21413, n21414, n21415, n21416, n21417, n21418, n21419, n21420,
         n21421, n21422, n21423, n21424, n21425, n21426, n21427, n21428,
         n21429, n21430, n21431, n21432, n21433, n21434, n21435, n21436,
         n21437, n21438, n21439, n21440, n21441, n21442, n21443, n21444,
         n21445, n21446, n21447, n21448, n21449, n21450, n21451, n21452,
         n21453, n21454, n21455, n21456, n21457, n21458, n21459, n21460,
         n21461, n21462, n21463, n21464, n21465, n21466, n21467, n21468,
         n21469, n21470, n21471, n21472, n21473, n21474, n21475, n21476,
         n21477, n21478, n21479, n21480, n21481, n21482, n21483, n21484,
         n21485, n21486, n21487, n21488, n21489, n21490, n21491, n21492,
         n21493, n21494, n21495, n21496, n21497, n21498, n21499, n21500,
         n21501, n21502, n21503, n21504, n21505, n21506, n21507, n21508,
         n21509, n21510, n21511, n21512, n21513, n21514, n21515, n21516,
         n21517, n21518, n21519, n21520, n21521, n21522, n21523, n21524,
         n21525, n21526, n21527, n21528, n21529, n21530, n21531, n21532,
         n21533, n21534, n21535, n21536, n21537, n21538, n21539, n21540,
         n21541, n21542, n21543, n21544, n21545, n21546, n21547, n21548,
         n21549, n21550, n21551, n21552, n21553, n21554, n21555, n21556,
         n21557, n21558, n21559, n21560, n21561, n21562, n21563, n21564,
         n21565, n21566, n21567, n21568, n21569, n21570, n21571, n21572,
         n21573, n21574, n21575, n21576, n21577, n21578, n21579, n21580,
         n21581, n21582, n21583, n21584, n21585, n21586, n21587, n21588,
         n21589, n21590, n21591, n21592, n21593, n21594, n21595, n21596,
         n21597, n21598, n21599, n21600, n21601, n21602, n21603, n21604,
         n21605, n21606, n21607, n21608, n21609, n21610, n21611, n21612,
         n21613, n21614, n21615, n21616, n21617, n21618, n21619, n21620,
         n21621, n21622, n21623, n21624, n21625, n21626, n21627, n21628,
         n21629, n21630, n21631, n21632, n21633, n21634, n21635, n21636,
         n21637, n21638, n21639, n21640, n21641, n21642, n21643, n21644,
         n21645, n21646, n21647, n21648, n21649, n21650, n21651, n21652,
         n21653, n21654, n21655, n21656, n21657, n21658, n21659, n21660,
         n21661, n21662, n21663, n21664, n21665, n21666, n21667, n21668,
         n21669, n21670, n21671, n21672, n21673, n21674, n21675, n21676,
         n21677, n21678, n21679, n21680, n21681, n21682, n21683, n21684,
         n21685, n21686, n21687, n21688, n21689, n21690, n21691, n21692,
         n21693, n21694, n21695, n21696, n21697, n21698, n21699, n21700,
         n21701, n21702, n21703, n21704, n21705, n21706, n21707, n21708,
         n21709, n21710, n21711, n21712, n21713, n21714, n21715, n21716,
         n21717, n21718, n21719, n21720, n21721, n21722, n21723, n21724,
         n21725, n21726, n21727, n21728, n21729, n21730, n21731, n21732,
         n21733, n21734, n21735, n21736, n21737, n21738, n21739, n21740,
         n21741, n21742, n21743, n21744, n21745, n21746, n21747, n21748,
         n21749, n21750, n21751, n21752, n21753, n21754, n21755, n21756,
         n21757, n21758, n21759, n21760, n21761, n21762, n21763, n21764,
         n21765, n21766, n21767, n21768, n21769, n21770, n21771, n21772,
         n21773, n21774, n21775, n21776, n21777, n21778, n21779, n21780,
         n21781, n21782, n21783, n21784, n21785, n21786, n21787, n21788,
         n21789, n21790, n21791, n21792, n21793, n21794, n21795, n21796,
         n21797, n21798, n21799, n21800, n21801, n21802, n21803, n21804,
         n21805, n21806, n21807, n21808, n21809, n21810, n21811, n21812,
         n21813, n21814, n21815, n21816, n21817, n21818, n21819, n21820,
         n21821, n21822, n21823, n21824, n21825, n21826, n21827, n21828,
         n21829, n21830, n21831, n21832, n21833, n21834, n21835, n21836,
         n21837, n21838, n21839, n21840, n21841, n21842, n21843, n21844,
         n21845, n21846, n21847, n21848, n21849, n21850, n21851, n21852,
         n21853, n21854, n21855, n21856, n21857, n21858, n21859, n21860,
         n21861, n21862, n21863, n21864, n21865, n21866, n21867, n21868,
         n21869, n21870, n21871, n21872, n21873, n21874, n21875, n21876,
         n21877, n21878, n21879, n21880, n21881, n21882, n21883, n21884,
         n21885, n21886, n21887, n21888, n21889, n21890, n21891, n21892,
         n21893, n21894, n21895, n21896, n21897, n21898, n21899, n21900,
         n21901, n21902, n21903, n21904, n21905, n21906, n21907, n21908,
         n21909, n21910, n21911, n21912, n21913, n21914, n21915, n21916,
         n21917, n21918, n21919, n21920, n21921, n21922, n21923, n21924,
         n21925, n21926, n21927, n21928, n21929, n21930, n21931, n21932,
         n21933, n21934, n21935, n21936, n21937, n21938, n21939, n21940,
         n21941, n21942, n21943, n21944, n21945, n21946, n21947, n21948,
         n21949, n21950, n21951, n21952, n21953, n21954, n21955, n21956,
         n21957, n21958, n21959, n21960, n21961, n21962, n21963, n21964,
         n21965, n21966, n21967, n21968, n21969, n21970, n21971, n21972,
         n21973, n21974, n21975, n21976, n21977, n21978, n21979, n21980,
         n21981, n21982, n21983, n21984, n21985, n21986, n21987, n21988,
         n21989, n21990, n21991, n21992, n21993, n21994, n21995, n21996,
         n21997, n21998, n21999, n22000, n22001, n22002, n22003, n22004,
         n22005, n22006, n22007, n22008, n22009, n22010, n22011, n22012,
         n22013, n22014, n22015, n22016, n22017, n22018, n22019, n22020,
         n22021, n22022, n22023, n22024, n22025, n22026, n22027, n22028,
         n22029, n22030, n22031, n22032, n22033, n22034, n22035, n22036,
         n22037, n22038, n22039, n22040, n22041, n22042, n22043, n22044,
         n22045, n22046, n22047, n22048, n22049, n22050, n22051, n22052,
         n22053, n22054, n22055, n22056, n22057, n22058, n22059, n22060,
         n22061, n22062, n22063, n22064, n22065, n22066, n22067, n22068,
         n22069, n22070, n22071, n22072, n22073, n22074, n22075, n22076,
         n22077, n22078, n22079, n22080, n22081, n22082, n22083, n22084,
         n22085, n22086, n22087, n22088, n22089, n22090, n22091, n22092,
         n22093, n22094, n22095, n22096, n22097, n22098, n22099, n22100,
         n22101, n22102, n22103, n22104, n22105, n22106, n22107, n22108,
         n22109, n22110, n22111, n22112, n22113, n22114, n22115, n22116,
         n22117, n22118, n22119, n22120, n22121, n22122, n22123, n22124,
         n22125, n22126, n22127, n22128, n22129, n22130, n22131, n22132,
         n22133, n22134, n22135, n22136, n22137, n22138, n22139, n22140,
         n22141, n22142, n22143, n22144, n22145, n22146, n22147, n22148,
         n22149, n22150, n22151, n22152, n22153, n22154, n22155, n22156,
         n22157, n22158, n22159, n22160, n22161, n22162, n22163, n22164,
         n22165, n22166, n22167, n22168, n22169, n22170, n22171, n22172,
         n22173, n22174, n22175, n22176, n22177, n22178, n22179, n22180,
         n22181, n22182, n22183, n22184, n22185, n22186, n22187, n22188,
         n22189, n22190, n22191, n22192, n22193, n22194, n22195, n22196,
         n22197, n22198, n22199, n22200, n22201, n22202, n22203, n22204,
         n22205, n22206, n22207, n22208, n22209, n22210, n22211, n22212,
         n22213, n22214, n22215, n22216, n22217, n22218, n22219, n22220,
         n22221, n22222, n22223, n22224, n22225, n22226, n22227, n22228,
         n22229, n22230, n22231, n22232, n22233, n22234, n22235, n22236,
         n22237, n22238, n22239, n22240, n22241, n22242, n22243, n22244,
         n22245, n22246, n22247, n22248, n22249, n22250, n22251, n22252,
         n22253, n22254, n22255, n22256, n22257, n22258, n22259, n22260,
         n22261, n22262, n22263, n22264, n22265, n22266, n22267, n22268,
         n22269, n22270, n22271, n22272, n22273, n22274, n22275, n22276,
         n22277, n22278, n22279, n22280, n22281, n22282, n22283, n22284,
         n22285, n22286, n22287, n22288, n22289, n22290, n22291, n22292,
         n22293, n22294, n22295, n22296, n22297, n22298, n22299, n22300,
         n22301, n22302, n22303, n22304, n22305, n22306, n22307, n22308,
         n22309, n22310, n22311, n22312, n22313, n22314, n22315, n22316,
         n22317, n22318, n22319, n22320, n22321, n22322, n22323, n22324,
         n22325, n22326, n22327, n22328, n22329, n22330, n22331, n22332,
         n22333, n22334, n22335, n22336, n22337, n22338, n22339, n22340,
         n22341, n22342, n22343, n22344, n22345, n22346, n22347, n22348,
         n22349, n22350, n22351, n22352, n22353, n22354, n22355, n22356,
         n22357, n22358, n22359, n22360, n22361, n22362, n22363, n22364,
         n22365, n22366, n22367, n22368, n22369, n22370, n22371, n22372,
         n22373, n22374, n22375, n22376, n22377, n22378, n22379, n22380,
         n22381, n22382, n22383, n22384, n22385, n22386, n22387, n22388,
         n22389, n22390, n22391, n22392, n22393, n22394, n22395, n22396,
         n22397, n22398, n22399, n22400, n22401, n22402, n22403, n22404,
         n22405, n22406, n22407, n22408, n22409, n22410, n22411, n22412,
         n22413, n22414, n22415, n22416, n22417, n22418, n22419, n22420,
         n22421, n22422, n22423, n22424, n22425, n22426, n22427, n22428,
         n22429, n22430, n22431, n22432, n22433, n22434, n22435, n22436,
         n22437, n22438, n22439, n22440, n22441, n22442, n22443, n22444,
         n22445, n22446, n22447, n22456, n22457, n22458, n22459, n22460,
         n22461, n22462, n22463, n22464, n22465, n22466, n22467, n22468,
         n22469, n22470, n22471, n22472, n22473, n22474, n22475, n22476,
         n22477, n22478, n22479, n22480, n22481, n22482, n22483, n22484,
         n22485, n22486, n22487, n22488, n22489, n22490, n22491, n22492,
         n22493, n22494, n22495, n22496, n22497, n22498, n22499, n22500,
         n22501, n22502, n22503, n22504, n22505, n22506, n22507, n22508,
         n22509, n22510, n22511, n22512, n22513, n22514, n22515, n22516,
         n22517, n22518, n22519, n22520, n22521, n22522, n22523, n22524,
         n22525, n22526, n22527, n22528, n22529, n22530, n22531, n22532,
         n22533, n22534, n22535, n22536, n22537, n22538, n22539, n22540,
         n22541, n22542, n22543, n22544, n22545, n22546, n22547, n22548,
         n22549, n22550, n22551, n22552, n22553, n22554, n22555, n22556,
         n22557, n22558, n22559, n22560, n22561, n22562, n22563, n22564,
         n22565, n22566, n22567, n22568, n22569, n22570, n22571, n22572,
         n22573, n22574, n22575, n22584, n22585, n22586, n22587, n22588,
         n22589, n22590, n22591, n22592, n22593, n22594, n22595, n22596,
         n22597, n22598, n22599, n22600, n22601, n22602, n22603, n22604,
         n22605, n22606, n22607, n22608, n22609, n22610, n22611, n22612,
         n22613, n22614, n22615, n22616, n22617, n22618, n22619, n22620,
         n22621, n22622, n22623, n22624, n22625, n22626, n22627, n22628,
         n22629, n22630, n22631, n22632, n22633, n22634, n22635, n22636,
         n22637, n22638, n22639, n22640, n22641, n22642, n22643, n22644,
         n22645, n22646, n22647, n22648, n22649, n22650, n22651, n22652,
         n22653, n22654, n22655, n22656, n22657, n22658, n22659, n22660,
         n22661, n22662, n22663, n22664, n22665, n22666, n22667, n22668,
         n22669, n22670, n22671, n22672, n22673, n22674, n22675, n22676,
         n22677, n22678, n22679, n22680, n22681, n22682, n22683, n22684,
         n22685, n22686, n22687, n22688, n22689, n22690, n22691, n22692,
         n22693, n22694, n22695, n22696, n22697, n22698, n22699, n22700,
         n22701, n22702, n22703, n22712, n22713, n22714, n22715, n22716,
         n22717, n22718, n22719, n22720, n22721, n22722, n22723, n22724,
         n22725, n22726, n22727, n22728, n22729, n22730, n22731, n22732,
         n22733, n22734, n22735, n22736, n22737, n22738, n22739, n22740,
         n22741, n22742, n22743, n22744, n22745, n22746, n22747, n22748,
         n22749, n22750, n22751, n22752, n22753, n22754, n22755, n22756,
         n22757, n22758, n22759, n22760, n22761, n22762, n22763, n22764,
         n22765, n22766, n22767, n22768, n22769, n22770, n22771, n22772,
         n22773, n22774, n22775, n22776, n22777, n22778, n22779, n22780,
         n22781, n22782, n22783, n22784, n22785, n22786, n22787, n22788,
         n22789, n22790, n22791, n22792, n22793, n22794, n22795, n22796,
         n22797, n22798, n22799, n22800, n22801, n22802, n22803, n22804,
         n22805, n22806, n22807, n22808, n22809, n22810, n22811, n22812,
         n22813, n22814, n22815, n22816, n22817, n22818, n22819, n22820,
         n22821, n22822, n22823, n22824, n22825, n22826, n22827, n22828,
         n22829, n22830, n22831, n22838, n22839, n22840, n22841, n22842,
         n22843, n22844, n22845, n22846, n22847, n22848, n22849, n22850,
         n22851, n22852, n22853, n22854, n22855, n22856, n22857, n22858,
         n22859, n22860, n22861, n22862, n22863, n22864, n22865, n22866,
         n22867, n22868, n22869, n22870, n22871, n22872, n22873, n22874,
         n22875, n22876, n22877, n22878, n22879, n22880, n22881, n22882,
         n22883, n22884, n22885, n22886, n22887, n22888, n22889, n22890,
         n22891, n22892, n22893, n22894, n22895, n22896, n22897, n22898,
         n22899, n22900, n22901, n22902, n22903, n22904, n22905, n22906,
         n22907, n22908, n22909, n22910, n22911, n22912, n22913, n22914,
         n22915, n22916, n22917, n22918, n22919, n22920, n22921, n22922,
         n22923, n22924, n22925, n22926, n22927, n22938, n22939, n22940,
         n22941, n22942, n22943, n22944, n22945, n22946, n22947, n22948,
         n22949, n22950, n22951, n22952, n22953, n22954, n22955, n22956,
         n22957, n22958, n22959, n22960, n22961, n22962, n22963, n22964,
         n22965, n22966, n22967, n22968, n22969, n22970, n22971, n22972,
         n22973, n22974, n22975, n22976, n22977, n22978, n22979, n22980,
         n22981, n22982, n22983, n22984, n22985, n22986, n22987, n22988,
         n22989, n22990, n22991, n22992, n22993, n22994, n22995, n22996,
         n22997, n22998, n22999, n23000, n23001, n23002, n23003, n23004,
         n23005, n23006, n23007, n23008, n23009, n23010, n23011, n23012,
         n23013, n23014, n23015, n23016, n23017, n23018, n23019, n23020,
         n23021, n23022, n23023, n23024, n23025, n23026, n23027, n23028,
         n23029, n23030, n23031, n23032, n23033, n23034, n23035, n23036,
         n23037, n23038, n23039, n23040, n23041, n23042, n23043, n23044,
         n23045, n23046, n23047, n23048, n23049, n23050, n23051, n23052,
         n23053, n23054, n23055, n23056, n23057, n23058, n23059, n23060,
         n23061, n23062, n23063, n23064, n23065, n23066, n23067, n23068,
         n23069, n23070, n23071, n23072, n23073, n23074, n23075, n23076,
         n23077, n23078, n23079, n23080, n23081, n23082, n23083, n23084,
         n23085, n23086, n23087, n23088, n23089, n23090, n23091, n23092,
         n23093, n23094, n23095, n23097, n23098, n23099, n23101, n23103,
         n23104, n23105, n23106, n23107, n23108, n23109, n23110, n23111,
         n23112, n23113, n23114, n23115, n23116, n23117, n23118, n23119,
         n23120, n23121, n23122, n23123, n23124, n23125, n23126, n23127,
         n23128, n23129, n23130, n23131, n23132, n23133, n23134, n23135,
         n23136, n23137, n23138, n23139, n23140, n23141, n23142, n23143,
         n23144, n23145, n23146, n23147, n23148, n23149, n23150, n23151,
         n23152, n23153, n23154, n23155, n23156, n23157, n23158, n23159,
         n23160, n23161, n23162, n23163, n23164, n23165, n23166, n23167,
         n23168, n23169, n23170, n23171, n23172, n23173, n23174, n23175,
         n23176, n23177, n23178, n23179, n23180, n23181, n23182, n23183,
         n23184, n23185, n23186, n23187, n23188, n23189, n23190, n23191,
         n23192, n23193, n23194, n23195, n23196, n23197, n23198, n23199,
         n23200, n23201, n23202, n23203, n23204, n23205, n23206, n23207,
         n23208, n23209, n23210, n23211, n23212, n23213, n23214, n23215,
         n23216, n23217, n23218, n23219, n23220, n23221, n23222, n23223,
         n23224, n23225, n23226, n23227, n23228, n23229, n23230, n23231,
         n23232, n23233, n23234, n23235, n23236, n23237, n23238, n23239,
         n23240, n23241, n23242, n23243, n23244, n23245, n23246, n23247,
         n23248, n23249, n23250, n23251, n23252, n23253, n23254, n23255,
         n23256, n23257, n23258, n23259, n23260, n23261, n23262, n23263,
         n23264, n23265, n23266, n23267, n23268, n23269, n23270, n23271,
         n23272, n23273, n23274, n23275, n23276, n23277, n23278, n23279,
         n23280, n23281, n23282, n23283, n23284, n23285, n23286, n23287,
         n23288, n23289, n23290, n23291, n23292, n23293, n23294, n23295,
         n23296, n23297, n23298, n23299, n23300, n23301, n23302, n23303,
         n23304, n23305, n23306, n23307, n23308, n23309, n23310, n23311,
         n23312, n23313, n23314, n23315, n23316, n23317, n23318, n23319,
         n23320, n23321, n23322, n23323, n23324, n23325, n23326, n23327,
         n23328, n23329, n23330, n23331, n23332, n23333, n23334, n23335,
         n23336, n23337, n23338, n23339, n23340, n23341, n23342, n23343,
         n23344, n23345, n23346, n23347, n23348, n23349, n23350, n23351,
         n23352, n23353, n23354, n23355, n23356, n23357, n23358, n23359,
         n23360, n23361, n23362, n23363, n23364, n23365, n23366, n23367,
         n23368, n23369, n23370, n23371, n23372, n23373, n23374, n23375,
         n23376, n23377, n23378, n23379, n23380, n23381, n23382, n23383,
         n23384, n23385, n23386, n23387, n23388, n23389, n23390, n23391,
         n23392, n23393, n23394, n23395, n23396, n23397, n23398, n23399,
         n23400, n23401, n23402, n23403, n23404, n23405, n23406, n23407,
         n23408, n23409, n23410, n23411, n23412, n23413, n23414, n23415,
         n23416, n23417, n23418, n23419, n23420, n23421, n23422, n23423,
         n23424, n23425, n23426, n23427, n23428, n23429, n23430, n23431,
         n23432, n23433, n23434, n23439, n23440, n23441, n23442, n23443,
         n23444, n23445, n23446, n23447, n23448, n23449, n23450, n23451,
         n23452, n23453, n23454, n23455, n23456, n23457, n23458, n23459,
         n23460, n23461, n23462, n23463, n23464, n23465, n23466, n23467,
         n23468, n23469, n23470, n23471, n23472, n23473, n23474, n23475,
         n23476, n23477, n23478, n23479, n23480, n23481, n23482, n23483,
         n23484, n23485, n23486, n23487, n23488, n23489, n23490, n23491,
         n23492, n23493, n23494, n23495, n23496, n23497, n23498, n23499,
         n23500, n23501, n23502, n23503, n23504, n23505, n23506, n23507,
         n23508, n23509, n23510, n23511, n23512, n23513, n23514, n23515,
         n23516, n23517, n23518, n23519, n23520, n23521, n23522, n23523,
         n23524, n23525, n23526, n23527, n23528, n23529, n23530, n23531,
         n23532, n23533, n23534, n23535, n23536, n23537, n23538, n23539,
         n23540, n23541, n23542, n23543, n23544, n23545, n23546, n23547,
         n23548, n23549, n23550, n23551, n23552, n23553, n23554, n23555,
         n23556, n23557, n23558, n23559, n23560, n23561, n23562, n23563,
         n23564, n23565, n23566, n23567, n23568, n23569, n23570, n23571,
         n23572, n23573, n23574, n23575, n23576, n23577, n23578, n23579,
         n23580, n23581, n23582, n23583, n23584, n23585, n23586, n23587,
         n23588, n23589, n23590, n23591, n23592, n23593, n23594, n23595,
         n23596, n23597, n23598, n23599, n23600, n23601, n23602, n23603,
         n23604, n23605, n23606, n23607, n23608, n23609, n23610, n23611,
         n23612, n23613, n23614, n23615, n23616, n23617, n23618, n23619,
         n23620, n23621, n23622, n23623, n23624, n23625, n23626, n23627,
         n23628, n23629, n23630, n23631, n23632, n23633, n23634, n23635,
         n23636, n23637, n23638, n23639, n23640, n23641, n23642, n23643,
         n23644, n23645, n23646, n23647, n23648, n23649, n23650, n23651,
         n23652, n23653, n23654, n23655, n23656, n23657, n23658, n23659,
         n23660, n23661, n23662, n23663, n23664, n23665, n23666, n23667,
         n23668, n23669, n23670, n23671, n23672, n23673, n23674, n23675,
         n23676, n23677, n23678, n23679, n23680, n23681, n23682, n23683,
         n23684, n23685, n23686, n23687, n23688, n23689, n23690, n23691,
         n23692, n23693, n23694, n23695, n23696, n23697, n23698, n23699,
         n23700, n23701, n23702, n23703, n23704, n23705, n23706, n23707,
         n23708, n23709, n23710, n23711, n23712, n23713, n23714, n23715,
         n23716, n23717, n23718, n23719, n23720, n23721, n23722, n23723,
         n23724, n23725, n23726, n23727, n23728, n23729, n23730, n23731,
         n23732, n23733, n23734, n23735, n23736, n23737, n23738, n23739,
         n23740, n23741, n23742, n23743, n23744, n23745, n23746, n23747,
         n23748, n23749, n23750, n23751, n23752, n23753, n23754, n23755,
         n23756, n23757, n23758, n23759, n23760, n23761, n23762, n23763,
         n23764, n23765, n23766, n23767, n23768, n23769, n23770, n23771,
         n23772, n23773, n23774, n23775, n23776, n23777, n23778, n23779,
         n23780, n23781, n23782, n23783, n23784, n23785, n23786, n23787,
         n23788, n23789, n23790, n23791, n23792, n23793, n23794, n23795,
         n23796, n23797, n23798, n23799, n23800, n23801, n23802, n23803,
         n23804, n23805, n23806, n23807, n23808, n23809, n23810, n23811,
         n23812, n23813, n23814, n23815, n23816, n23817, n23818, n23819,
         n23820, n23821, n23822, n23823, n23824, n23825, n23826, n23827,
         n23828, n23829, n23830, n23831, n23832, n23833, n23834, n23835,
         n23836, n23837, n23838, n23839, n23840, n23841, n23842, n23843,
         n23844, n23845, n23846, n23847, n23848, n23849, n23850, n23851,
         n23852, n23853, n23854, n23855, n23856, n23857, n23858, n23859,
         n23860, n23861, n23862, n23863, n23864, n23865, n23866, n23867,
         n23868, n23869, n23870, n23871, n23872, n23873, n23874, n23875,
         n23876, n23877, n23878, n23879, n23880, n23881, n23882, n23883,
         n23884, n23885, n23886, n23887, n23888, n23889, n23890, n23891,
         n23892, n23893, n23894, n23895, n23896, n23897, n23898, n23899,
         n23900, n23901, n23902, n23903, n23904, n23905, n23906, n23907,
         n23908, n23909, n23910, n23911, n23912, n23913, n23914, n23915,
         n23916, n23917, n23918, n23919, n23920, n23921, n23922, n23923,
         n23924, n23925, n23926, n23927, n23928, n23929, n23930, n23931,
         n23932, n23933, n23934, n23935, n23936, n23937, n23938, n23939,
         n23940, n23941, n23942, n23943, n23944, n23945, n23946, n23947,
         n23948, n23949, n23950, n23951, n23952, n23953, n23954, n23955,
         n23956, n23957, n23958, n23959, n23960, n23961, n23962, n23963,
         n23964, n23965, n23966, n23967, n23968, n23969, n23970, n23971,
         n23972, n23973, n23974, n23975, n23976, n23977, n23978, n23979,
         n23980, n23981, n23982, n23983, n23984, n23985, n23986, n23987,
         n23988, n23989, n23990, n23991, n23992, n23993, n23994, n23995,
         n23996, n23997, n23998, n23999, n24000, n24001, n24002, n24003,
         n24004, n24005, n24006, n24007, n24008, n24009, n24010, n24011,
         n24012, n24013, n24014, n24015, n24016, n24017, n24018, n24019,
         n24020, n24021, n24022, n24023, n24024, n24025, n24026, n24027,
         n24028, n24029, n24030, n24031, n24032, n24033, n24034, n24035,
         n24036, n24037, n24038, n24039, n24040, n24041, n24042, n24043,
         n24044, n24045, n24046, n24047, n24048, n24049, n24050, n24051,
         n24052, n24053, n24054, n24055, n24056, n24057, n24058, n24059,
         n24060, n24061, n24062, n24063, n24064, n24065, n24066, n24067,
         n24068, n24069, n24070, n24071, n24072, n24073, n24074, n24075,
         n24076, n24077, n24078, n24079, n24080, n24081, n24082, n24083,
         n24084, n24085, n24086, n24087, n24088, n24089, n24090, n24091,
         n24092, n24093, n24094, n24095, n24096, n24097, n24098, n24099,
         n24100, n24101, n24102, n24103, n24104, n24105, n24106, n24107,
         n24108, n24109, n24110, n24111, n24112, n24113, n24114, n24115,
         n24116, n24117, n24118, n24119, n24120, n24121, n24122, n24123,
         n24124, n24125, n24126, n24127, n24128, n24129, n24130, n24131,
         n24132, n24133, n24134, n24135, n24136, n24137, n24138, n24139,
         n24140, n24141, n24142, n24143, n24144, n24145, n24146, n24147,
         n24148, n24149, n24150, n24151, n24152, n24153, n24154, n24155,
         n24156, n24157, n24158, n24159, n24160, n24161, n24162, n24163,
         n24164, n24165, n24166, n24167, n24168, n24169, n24170, n24171,
         n24172, n24173, n24174, n24175, n24176, n24177, n24178, n24179,
         n24180, n24181, n24182, n24183, n24184, n24185, n24186, n24187,
         n24188, n24189, n24190, n24191, n24192, n24193, n24194, n24195,
         n24196, n24197, n24198, n24199, n24200, n24201, n24202, n24203,
         n24204, n24205, n24206, n24207, n24208, n24209, n24210, n24211,
         n24212, n24213, n24214, n24215, n24216, n24217, n24218, n24219,
         n24220, n24221, n24222, n24223, n24224, n24225, n24226, n24227,
         n24228, n24229, n24230, n24231, n24232, n24233, n24234, n24235,
         n24236, n24237, n24238, n24239, n24240, n24241, n24242, n24243,
         n24244, n24245, n24246, n24247, n24248, n24249, n24250, n24251,
         n24252, n24253, n24254, n24255, n24256, n24257, n24258, n24259,
         n24260, n24261, n24262, n24263, n24264, n24265, n24266, n24267,
         n24268, n24269, n24270, n24271, n24272, n24273, n24274, n24275,
         n24276, n24277, n24278, n24279, n24280, n24281, n24282, n24283,
         n24284, n24285, n24286, n24287, n24288, n24289, n24290, n24291,
         n24292, n24293, n24294, n24295, n24296, n24297, n24298, n24299,
         n24300, n24301, n24302, n24303, n24304, n24305, n24306, n24307,
         n24308, n24309, n24310, n24311, n24312, n24313, n24314, n24315,
         n24316, n24317, n24318, n24319, n24320, n24321, n24322, n24323,
         n24324, n24325, n24326, n24327, n24328, n24329, n24330, n24331,
         n24332, n24333, n24334, n24335, n24336, n24337, n24338, n24339,
         n24340, n24341, n24342, n24343, n24344, n24345, n24346, n24347,
         n24348, n24349, n24350, n24351, n24352, n24353, n24354, n24355,
         n24356, n24357, n24358, n24359, n24360, n24361, n24362, n24363,
         n24364, n24365, n24366, n24367, n24368, n24369, n24370, n24371,
         n24372, n24373, n24374, n24375, n24376, n24377, n24378, n24379,
         n24380, n24381, n24382, n24383, n24384, n24385, n24386, n24387,
         n24388, n24389, n24390, n24391, n24392, n24393, n24394, n24395,
         n24396, n24397, n24398, n24399, n24400, n24401, n24402, n24403,
         n24404, n24405, n24406, n24407, n24408, n24409, n24410, n24411,
         n24412, n24413, n24414, n24415, n24416, n24417, n24418, n24419,
         n24420, n24421, n24422, n24423, n24424, n24425, n24426, n24427,
         n24428, n24429, n24430, n24431, n24432, n24433, n24434, n24435,
         n24436, n24437, n24438, n24439, n24440, n24441, n24442, n24443,
         n24444, n24445, n24446, n24447, n24448, n24449, n24450, n24451,
         n24452, n24453, n24454, n24455, n24456, n24457, n24458, n24459,
         n24460, n24461, n24462, n24463, n24464, n24465, n24466, n24467,
         n24468, n24469, n24470, n24471, n24472, n24473, n24474, n24475,
         n24476, n24477, n24478, n24479, n24480, n24481, n24482, n24483,
         n24484, n24485, n24486, n24487, n24488, n24489, n24490, n24491,
         n24492, n24493, n24494, n24495, n24496, n24497, n24498, n24499,
         n24500, n24501, n24502, n24503, n24504, n24505, n24506, n24507,
         n24508, n24509, n24510, n24511, n24512, n24513, n24514, n24515,
         n24516, n24517, n24518, n24519, n24520, n24521, n24522, n24523,
         n24524, n24525, n24526, n24527, n24528, n24529, n24530, n24531,
         n24532, n24533, n24534, n24535, n24536, n24537, n24538, n24539,
         n24540, n24541, n24542, n24543, n24544, n24545, n24546, n24547,
         n24548, n24549, n24550, n24551, n24552, n24553, n24554, n24555,
         n24556, n24557, n24558, n24559, n24560, n24561, n24562, n24563,
         n24564, n24565, n24566, n24567, n24568, n24569, n24570, n24571,
         n24572, n24573, n24574, n24575, n24576, n24577, n24578, n24579,
         n24580, n24581, n24582, n24583, n24584, n24585, n24586, n24587,
         n24588, n24589, n24590, n24591, n24592, n24593, n24594, n24595,
         n24596, n24597, n24598, n24599, n24600, n24601, n24602, n24603,
         n24604, n24605, n24606, n24607, n24608, n24609, n24610, n24611,
         n24612, n24613, n24614, n24615, n24616, n24617, n24618, n24619,
         n24620, n24621, n24622, n24623, n24624, n24625, n24626, n24627,
         n24628, n24629, n24630, n24631, n24632, n24633, n24634, n24635,
         n24636, n24637, n24638, n24639, n24640, n24641, n24642, n24643,
         n24644, n24645, n24646, n24647, n24648, n24649, n24650, n24651,
         n24652, n24653, n24654, n24655, n24656, n24657, n24658, n24659,
         n24660, n24661, n24662, n24663, n24664, n24665, n24666, n24667,
         n24668, n24669, n24670, n24671, n24672, n24673, n24674, n24675,
         n24676, n24677, n24678, n24679, n24680, n24681, n24682, n24683,
         n24684, n24685, n24686, n24687, n24688, n24689, n24690, n24691,
         n24692, n24693, n24694, n24695, n24696, n24697, n24698, n24699,
         n24700, n24701, n24702, n24703, n24704, n24705, n24706, n24707,
         n24708, n24709, n24710, n24711, n24712, n24713, n24714, n24715,
         n24716, n24717, n24718, n24719, n24720, n24721, n24722, n24723,
         n24724, n24725, n24726, n24727, n24728, n24729, n24730, n24731,
         n24732, n24733, n24734, n24735, n24736, n24737, n24738, n24739,
         n24740, n24741, n24742, n24743, n24744, n24745, n24746, n24747,
         n24748, n24749, n24750, n24751, n24752, n24753, n24754, n24755,
         n24756, n24757, n24758, n24759, n24760, n24761, n24762, n24763,
         n24764, n24765, n24766, n24767, n24768, n24769, n24770, n24771,
         n24772, n24773, n24774, n24775, n24776, n24777, n24778, n24779,
         n24780, n24781, n24782, n24783, n24784, n24785, n24786, n24787,
         n24788, n24789, n24790, n24791, n24792, n24793, n24794, n24795,
         n24796, n24797, n24798, n24799, n24800, n24801, n24802, n24803,
         n24804, n24805, n24806, n24807, n24808, n24809, n24810, n24811,
         n24812, n24813, n24814, n24815, n24816, n24817, n24818, n24819,
         n24820, n24821, n24822, n24823, n24832, n24833, n24834, n24835,
         n24836, n24837, n24838, n24839, n24840, n24841, n24842, n24843,
         n24844, n24845, n24846, n24847, n24848, n24849, n24850, n24851,
         n24852, n24853, n24854, n24855, n24856, n24857, n24858, n24859,
         n24860, n24861, n24862, n24863, n24864, n24865, n24866, n24867,
         n24868, n24869, n24870, n24871, n24872, n24873, n24874, n24875,
         n24876, n24877, n24878, n24879, n24880, n24881, n24882, n24883,
         n24884, n24885, n24886, n24887, n24888, n24889, n24890, n24891,
         n24892, n24893, n24894, n24895, n24896, n24897, n24898, n24899,
         n24900, n24901, n24902, n24903, n24904, n24905, n24906, n24907,
         n24908, n24909, n24910, n24911, n24912, n24913, n24914, n24915,
         n24916, n24917, n24918, n24919, n24920, n24921, n24922, n24923,
         n24924, n24925, n24926, n24927, n24928, n24929, n24930, n24931,
         n24932, n24933, n24934, n24935, n24936, n24937, n24938, n24939,
         n24940, n24941, n24942, n24943, n24944, n24945, n24946, n24947,
         n24948, n24949, n24950, n24951, n24952, n24953, n24954, n24955,
         n24956, n24957, n24958, n24959, n24960, n24961, n24962, n24963,
         n24964, n24965, n24966, n24967, n24968, n24969, n24970, n24971,
         n24972, n24973, n24974, n24975, n24976, n24977, n24978, n24979,
         n24980, n24981, n24982, n24983, n24984, n24985, n24986, n24987,
         n24988, n24989, n24990, n24991, n24992, n24993, n24994, n24995,
         n24996, n24997, n24998, n24999, n25000, n25001, n25002, n25003,
         n25004, n25005, n25006, n25007, n25008, n25009, n25010, n25011,
         n25012, n25013, n25014, n25015, n25016, n25017, n25018, n25019,
         n25020, n25021, n25022, n25023, n25024, n25025, n25026, n25027,
         n25028, n25029, n25030, n25031, n25032, n25033, n25034, n25035,
         n25036, n25037, n25038, n25039, n25040, n25041, n25042, n25043,
         n25044, n25045, n25046, n25047, n25048, n25049, n25050, n25051,
         n25052, n25053, n25054, n25055, n25056, n25057, n25058, n25059,
         n25060, n25061, n25062, n25063, n25064, n25065, n25066, n25067,
         n25068, n25069, n25070, n25071, n25072, n25073, n25074, n25075,
         n25076, n25077, n25078, n25079, n25080, n25081, n25082, n25083,
         n25084, n25085, n25086, n25087, n25088, n25089, n25090, n25091,
         n25092, n25093, n25094, n25095, n25096, n25097, n25098, n25099,
         n25100, n25101, n25102, n25103, n25104, n25105, n25106, n25107,
         n25108, n25109, n25110, n25111, n25112, n25113, n25114, n25115,
         n25116, n25117, n25118, n25119, n25120, n25121, n25122, n25123,
         n25124, n25125, n25126, n25127, n25128, n25129, n25130, n25131,
         n25132, n25133, n25134, n25135, n25136, n25137, n25138, n25139,
         n25140, n25141, n25142, n25143, n25144, n25145, n25146, n25147,
         n25148, n25149, n25150, n25151, n25152, n25153, n25154, n25155,
         n25156, n25157, n25158, n25159, n25160, n25161, n25162, n25163,
         n25164, n25165, n25166, n25167, n25168, n25169, n25170, n25171,
         n25172, n25173, n25174, n25175, n25176, n25177, n25178, n25179,
         n25180, n25181, n25182, n25183, n25184, n25185, n25186, n25187,
         n25188, n25189, n25190, n25191, n25192, n25193, n25194, n25195,
         n25196, n25197, n25198, n25199, n25200, n25201, n25202, n25203,
         n25204, n25205, n25206, n25207, n25208, n25209, n25210, n25211,
         n25212, n25213, n25214, n25215, n25216, n25217, n25218, n25219,
         n25220, n25221, n25222, n25223, n25224, n25225, n25226, n25227,
         n25228, n25229, n25230, n25231, n25232, n25233, n25234, n25235,
         n25236, n25237, n25238, n25239, n25240, n25241, n25242, n25243,
         n25244, n25245, n25246, n25247, n25248, n25249, n25250, n25251,
         n25252, n25253, n25254, n25255, n25256, n25257, n25258, n25259,
         n25260, n25261, n25262, n25263, n25264, n25265, n25266, n25267,
         n25268, n25269, n25270, n25271, n25272, n25273, n25274, n25275,
         n25276, n25277, n25278, n25279, n25280, n25281, n25282, n25283,
         n25284, n25285, n25286, n25287, n25288, n25289, n25290, n25291,
         n25292, n25293, n25294, n25295, n25296, n25297, n25298, n25299,
         n25300, n25301, n25302, n25303, n25304, n25305, n25306, n25307,
         n25308, n25309, n25310, n25311, n25312, n25313, n25314, n25315,
         n25316, n25317, n25318, n25319, n25320, n25321, n25322, n25323,
         n25324, n25325, n25326, n25327, n25328, n25329, n25330, n25331,
         n25332, n25333, n25334, n25335, n25336, n25337, n25338, n25339,
         n25340, n25341, n25342, n25343, n25344, n25345, n25346, n25347,
         n25348, n25349, n25350, n25351, n25352, n25353, n25354, n25355,
         n25356, n25357, n25358, n25359, n25360, n25361, n25362, n25363,
         n25364, n25365, n25366, n25367, n25368, n25369, n25370, n25371,
         n25372, n25373, n25374, n25375, n25376, n25377, n25378, n25379,
         n25380, n25381, n25382, n25383, n25384, n25385, n25386, n25387,
         n25388, n25389, n25390, n25391, n25392, n25393, n25394, n25395,
         n25396, n25397, n25398, n25399, n25400, n25401, n25402, n25403,
         n25404, n25405, n25406, n25407, n25408, n25409, n25410, n25411,
         n25412, n25413, n25414, n25415, n25416, n25417, n25418, n25419,
         n25420, n25421, n25422, n25423, n25424, n25425, n25426, n25427,
         n25428, n25429, n25430, n25431, n25432, n25433, n25434, n25435,
         n25436, n25437, n25438, n25439, n25440, n25441, n25442, n25443,
         n25444, n25445, n25446, n25447, n25448, n25449, n25450, n25451,
         n25452, n25453, n25454, n25455, n25456, n25457, n25458, n25459,
         n25460, n25461, n25462, n25463, n25464, n25465, n25466, n25467,
         n25468, n25469, n25470, n25471, n25472, n25473, n25474, n25475,
         n25476, n25477, n25478, n25479, n25480, n25481, n25482, n25483,
         n25484, n25485, n25486, n25487, n25488, n25489, n25490, n25491,
         n25492, n25493, n25494, n25495, n25496, n25497, n25498, n25499,
         n25500, n25501, n25502, n25503, n25504, n25505, n25506, n25507,
         n25508, n25509, n25510, n25511, n25512, n25513, n25514, n25515,
         n25516, n25517, n25518, n25519, n25520, n25521, n25522, n25523,
         n25524, n25525, n25526, n25527, n25528, n25529, n25530, n25531,
         n25532, n25533, n25534, n25535, n25536, n25537, n25538, n25539,
         n25540, n25541, n25542, n25543, n25544, n25545, n25546, n25547,
         n25548, n25549, n25550, n25551, n25552, n25553, n25554, n25555,
         n25556, n25557, n25558, n25559, n25560, n25561, n25562, n25563,
         n25564, n25565, n25566, n25567, n25568, n25569, n25570, n25571,
         n25572, n25573, n25574, n25575, n25576, n25577, n25578, n25579,
         n25580, n25581, n25582, n25583, n25584, n25585, n25586, n25587,
         n25588, n25589, n25590, n25591, n25592, n25593, n25594, n25595,
         n25596, n25597, n25598, n25599, n25600, n25601, n25602, n25603,
         n25604, n25605, n25606, n25607, n25608, n25609, n25610, n25611,
         n25612, n25613, n25614, n25615, n25616, n25617, n25618, n25619,
         n25620, n25621, n25622, n25623, n25624, n25625, n25626, n25627,
         n25628, n25629, n25630, n25631, n25632, n25633, n25634, n25635,
         n25636, n25637, n25638, n25639, n25640, n25641, n25642, n25643,
         n25644, n25645, n25646, n25647, n25648, n25649, n25650, n25651,
         n25652, n25653, n25654, n25655, n25656, n25657, n25658, n25659,
         n25660, n25661, n25662, n25663, n25664, n25665, n25666, n25667,
         n25668, n25669, n25670, n25671, n25672, n25673, n25674, n25675,
         n25676, n25677, n25678, n25679, n25680, n25681, n25682, n25683,
         n25684, n25685, n25686, n25687, n25688, n25689, n25690, n25691,
         n25692, n25693, n25694, n25695, n25696, n25697, n25698, n25699,
         n25700, n25701, n25702, n25703, n25704, n25705, n25706, n25707,
         n25708, n25709, n25710, n25711, n25712, n25713, n25714, n25715,
         n25716, n25717, n25718, n25719, n25720, n25721, n25722, n25723,
         n25724, n25725, n25726, n25727, n25728, n25729, n25730, n25731,
         n25732, n25735, n25736, n25737, n25738, n25739, n25740, n25741,
         n25742, n25743, n25744, n25745, n25746, n25747, n25748, n25749,
         n25750, n25751, n25752, n25753, n25754, n25755, n25756, n25757,
         n25758, n25759, n25760, n25761, n25762, n25763, n25764, n25765,
         n25766, n25767, n25768, n25769, n25770, n25771, n25772, n25773,
         n25774, n25775, n25776, n25777, n25778, n25779, n25780, n25781,
         n25782, n25783, n25784, n25785, n25786, n25787, n25788, n25789,
         n25790, n25791, n25792, n25793, n25794, n25795, n25796, n25797,
         n25798, n25799, n25800, n25801, n25802, n25803, n25804, n25805,
         n25806, n25807, n25808, n25809, n25810, n25811, n25812, n25813,
         n25814, n25815, n25816, n25817, n25818, n25819, n25820, n25821,
         n25822, n25823, n25824, n25825, n25826, n25827, n25828, n25829,
         n25830, n25831, n25832, n25833, n25834, n25835, n25836, n25837,
         n25838, n25839, n25840, n25841, n25842, n25843, n25844, n25845,
         n25846, n25847, n25848, n25849, n25850, n25851, n25852, n25853,
         n25854, n25855, n25856, n25857, n25858, n25859, n25860, n25861,
         n25862, n25863, n25864, n25865, n25866, n25867, n25868, n25869,
         n25870, n25871, n25872, n25873, n25874, n25875, n25876, n25877,
         n25878, n25879, n25880, n25881, n25882, n25883, n25884, n25885,
         n25886, n25887, n25888, n25889, n25890, n25891, n25892, n25893,
         n25894, n25895, n25896, n25897, n25898, n25899, n25900, n25901,
         n25902, n25903, n25904, n25905, n25906, n25907, n25908, n25909,
         n25910, n25911, n25912, n25913, n25914, n25915, n25916, n25917,
         n25918, n25919, n25920, n25921, n25922, n25923, n25924, n25925,
         n25926, n25927, n25928, n25929, n25930, n25931, n25932, n25933,
         n25934, n25935, n25936, n25937, n25938, n25939, n25940, n25941,
         n25942, n25943, n25944, n25945, n25946, n25947, n25948, n25949,
         n25950, n25951, n25952, n25953, n25954, n25955, n25956, n25957,
         n25958, n25959, n25960, n25961, n25962, n25963, n25964, n25965,
         n25966, n25967, n25968, n25969, n25970, n25971, n25972, n25973,
         n25974, n25975, n25976, n25977, n25978, n25979, n25980, n25981,
         n25982, n25983, n25984, n25985, n25986, n25987, n25988, n25989,
         n25990, n25991, n25992, n25993, n25994, n25995, n25996, n25997,
         n25998, n25999, n26000, n26001, n26002, n26003, n26004, n26005,
         n26006, n26007, n26008, n26009, n26010, n26011, n26012, n26013,
         n26014, n26015, n26016, n26017, n26018, n26019, n26020, n26021,
         n26022, n26023, n26024, n26025, n26026, n26027, n26028, n26029,
         n26030, n26031, n26032, n26033, n26034, n26035, n26036, n26037,
         n26038, n26039, n26040, n26041, n26042, n26043, n26044, n26045,
         n26046, n26047, n26048, n26049, n26050, n26051, n26052, n26053,
         n26054, n26055, n26056, n26057, n26058, n26059, n26060, n26061,
         n26062, n26063, n26064, n26065, n26066, n26067, n26068, n26069,
         n26070, n26071, n26072, n26073, n26074, n26075, n26076, n26077,
         n26078, n26079, n26080, n26081, n26082, n26083, n26084, n26085,
         n26086, n26087, n26088, n26089, n26090, n26091, n26092, n26093,
         n26094, n26095, n26096, n26097, n26098, n26099, n26100, n26101,
         n26102, n26103, n26104, n26105, n26106, n26107, n26108, n26109,
         n26110, n26111, n26112, n26113, n26114, n26115, n26116, n26117,
         n26118, n26119, n26120, n26121, n26122, n26123, n26124, n26125,
         n26126, n26127, n26128, n26129, n26130, n26131, n26132, n26133,
         n26134, n26135, n26136, n26137, n26138, n26139, n26140, n26141,
         n26142, n26143, n26144, n26145, n26146, n26147, n26148, n26149,
         n26150, n26151, n26152, n26153, n26154, n26155, n26156, n26157,
         n26158, n26159, n26160, n26161, n26162, n26163, n26164, n26165,
         n26166, n26167, n26168, n26169, n26170, n26171, n26172, n26173,
         n26174, n26175, n26176, n26177, n26178, n26179, n26180, n26181,
         n26182, n26183, n26184, n26185, n26186, n26187, n26188, n26189,
         n26190, n26191, n26192, n26193, n26194, n26195, n26196, n26197,
         n26198, n26199, n26200, n26201, n26202, n26203, n26204, n26205,
         n26206, n26207, n26208, n26209, n26210, n26211, n26212, n26213,
         n26214, n26215, n26216, n26217, n26218, n26219, n26220, n26221,
         n26222, n26223, n26224, n26225, n26226, n26227, n26228, n26229,
         n26230, n26231, n26232, n26233, n26234, n26235, n26236, n26237,
         n26238, n26239, n26240, n26241, n26242, n26243, n26244, n26245,
         n26246, n26247, n26248, n26249, n26250, n26251, n26252, n26253,
         n26254, n26255, n26256, n26257, n26258, n26259, n26260, n26261,
         n26262, n26263, n26264, n26265, n26266, n26267, n26268, n26269,
         n26270, n26271, n26272, n26273, n26274, n26275, n26276, n26277,
         n26278, n26279, n26280, n26281, n26282, n26283, n26284, n26285,
         n26286, n26287, n26288, n26289, n26290, n26291, n26292, n26293,
         n26294, n26295, n26296, n26297, n26298, n26299, n26300, n26301,
         n26302, n26303, n26304, n26305, n26306, n26307, n26308, n26309,
         n26310, n26311, n26312, n26313, n26314, n26315, n26316, n26317,
         n26318, n26319, n26320, n26321, n26322, n26323, n26324, n26325,
         n26326, n26327, n26328, n26329, n26330, n26331, n26332, n26333,
         n26334, n26335, n26336, n26337, n26338, n26339, n26340, n26341,
         n26342, n26343, n26344, n26345, n26346, n26347, n26348, n26349,
         n26350, n26351, n26352, n26353, n26354, n26355, n26356, n26357,
         n26358, n26359, n26360, n26361, n26362, n26363, n26364, n26365,
         n26366, n26367, n26368, n26369, n26370, n26371, n26372, n26373,
         n26374, n26375, n26376, n26377, n26378, n26379, n26380, n26381,
         n26382, n26383, n26384, n26385, n26386, n26387, n26388, n26389,
         n26390, n26391, n26392, n26393, n26394, n26395, n26396, n26397,
         n26398, n26399, n26400, n26401, n26402, n26403, n26404, n26405,
         n26406, n26407, n26408, n26409, n26410, n26411, n26412, n26413,
         n26414, n26415, n26416, n26417, n26418, n26419, n26420, n26421,
         n26422, n26423, n26424, n26425, n26426, n26427, n26428, n26429,
         n26430, n26431, n26432, n26433, n26434, n26435, n26436, n26437,
         n26438, n26439, n26440, n26441, n26442, n26443, n26444, n26445,
         n26446, n26447, n26448, n26449, n26450, n26451, n26452, n26453,
         n26454, n26455, n26456, n26457, n26458, n26459, n26460, n26461,
         n26462, n26463, n26464, n26465, n26466, n26467, n26468, n26469,
         n26470, n26471, n26472, n26473, n26474, n26475, n26476, n26477,
         n26478, n26479, n26480, n26481, n26482, n26483, n26484, n26485,
         n26486, n26487, n26488, n26489, n26490, n26491, n26492, n26493,
         n26494, n26495, n26496, n26497, n26498, n26499, n26500, n26501,
         n26502, n26503, n26504, n26505, n26506, n26507, n26508, n26509,
         n26510, n26511, n26512, n26513, n26514, n26515, n26516, n26517,
         n26518, n26519, n26520, n26521, n26522, n26523, n26524, n26525,
         n26526, n26527, n26528, n26529, n26530, n26531, n26532, n26533,
         n26534, n26535, n26536, n26537, n26538, n26539, n26540, n26541,
         n26542, n26543, n26544, n26545, n26546, n26547, n26548, n26549,
         n26550, n26551, n26552, n26553, n26554, n26555, n26556, n26557,
         n26558, n26559, n26560, n26561, n26562, n26563, n26564, n26565,
         n26566, n26567, n26568, n26569, n26570, n26571, n26572, n26573,
         n26574, n26575, n26576, n26577, n26578, n26579, n26580, n26581,
         n26582, n26583, n26584, n26585, n26586, n26587, n26588, n26589,
         n26590, n26591, n26592, n26593, n26594, n26595, n26596, n26597,
         n26598, n26599, n26600, n26601, n26602, n26603, n26604, n26605,
         n26606, n26607, n26608, n26609, n26610, n26611, n26612, n26613,
         n26614, n26615, n26616, n26617, n26618, n26619, n26620, n26621,
         n26622, n26623, n26624, n26625, n26626, n26627, n26628, n26629,
         n26630, n26631, n26632, n26633, n26634, n26635, n26636, n26637,
         n26638, n26639, n26640, n26641, n26642, n26643, n26644, n26645,
         n26646, n26647, n26648, n26649, n26650, n26651, n26652, n26653,
         n26654, n26655, n26656, n26657, n26658, n26659, n26660, n26661,
         n26662, n26663, n26664, n26665, n26666, n26667, n26668, n26669,
         n26670, n26671, n26672, n26673, n26674, n26675, n26676, n26677,
         n26678, n26679, n26680, n26681, n26682, n26683, n26684, n26685,
         n26686, n26687, n26688, n26689, n26690, n26691, n26692, n26693,
         n26694, n26695, n26696, n26697, n26698, n26699, n26700, n26701,
         n26702, n26703, n26704, n26705, n26706, n26707, n26708, n26709,
         n26710, n26711, n26712, n26713, n26714, n26715, n26716, n26717,
         n26718, n26719, n26720, n26721, n26722, n26723, n26724, n26725,
         n26726, n26727, n26728, n26729, n26730, n26731, n26732, n26733,
         n26734, n26735, n26736, n26737, n26738, n26739, n26740, n26741,
         n26742, n26743, n26744, n26745, n26746, n26747, n26748, n26749,
         n26750, n26751, n26752, n26753, n26754, n26755, n26756, n26757,
         n26758, n26759, n26760, n26761, n26762, n26763, n26764, n26765,
         n26766, n26767, n26768, n26769, n26770, n26771, n26772, n26773,
         n26774, n26775, n26776, n26777, n26778, n26779, n26780, n26781,
         n26782, n26783, n26784, n26785, n26786, n26787, n26788, n26789,
         n26790, n26791, n26792, n26793, n26794, n26795, n26796, n26797,
         n26798, n26799, n26800, n26801, n26802, n26803, n26804, n26805,
         n26806, n26807, n26808, n26809, n26810, n26811, n26812, n26813,
         n26814, n26815, n26816, n26817, n26818, n26819, n26820, n26821,
         n26822, n26823, n26824, n26825, n26826, n26827, n26828, n26829,
         n26830, n26831, n26832, n26833, n26834, n26835, n26836, n26837,
         n26838, n26839, n26840, n26841, n26842, n26843, n26844, n26845,
         n26846, n26847, n26848, n26849, n26850, n26851, n26852, n26853,
         n26854, n26855, n26856, n26857, n26858, n26859, n26860, n26861,
         n26862, n26863, n26864, n26865, n26866, n26867, n26868, n26869,
         n26870, n26871, n26872, n26873, n26874, n26875, n26876, n26877,
         n26878, n26879, n26880, n26881, n26882, n26883, n26884, n26885,
         n26886, n26887, n26888, n26889, n26890, n26891, n26892, n26893,
         n26894, n26895, n26896, n26897, n26898, n26899, n26900, n26901,
         n26902, n26903, n26904, n26905, n26906, n26907, n26908, n26909,
         n26910, n26911, n26912, n26913, n26914, n26915, n26916, n26917,
         n26918, n26919, n26920, n26921, n26922, n26923, n26924, n26925,
         n26926, n26927, n26928, n26929, n26930, n26931, n26932, n26933,
         n26934, n26935, n26936, n26937, n26938, n26939, n26940, n26941,
         n26942, n26943, n26944, n26945, n26946, n26947, n26948, n26949,
         n26950, n26951, n26952, n26953, n26954, n26955, n26956, n26957,
         n26958, n26959, n26960, n26961, n26962, n26963, n26964, n26965,
         n26966, n26967, n26968, n26969, n26970, n26971, n26972, n26973,
         n26974, n26975, n26976, n26977, n26978, n26979, n26980, n26981,
         n26982, n26983, n26984, n26985, n26986, n26987, n26988, n26989,
         n26990, n26991, n26992, n26993, n26994, n26995, n26996, n26997,
         n26998, n26999, n27000, n27001, n27002, n27003, n27004, n27005,
         n27006, n27007, n27008, n27009, n27010, n27011, n27012, n27013,
         n27014, n27015, n27016, n27017, n27018, n27019, n27020, n27021,
         n27022, n27023, n27024, n27025, n27026, n27027, n27028, n27029,
         n27030, n27031, n27032, n27033, n27034, n27035, n27036, n27037,
         n27038, n27039, n27040, n27041, n27042, n27043, n27044, n27045,
         n27046, n27047, n27048, n27049, n27050, n27051, n27052, n27053,
         n27054, n27055, n27056, n27057, n27058, n27059, n27060, n27061,
         n27062, n27063, n27064, n27065, n27066, n27067, n27068, n27069,
         n27070, n27071, n27072, n27073, n27074, n27075, n27076, n27077,
         n27078, n27079, n27080, n27081, n27082, n27083, n27084, n27085,
         n27086, n27087, n27088, n27089, n27090, n27091, n27092, n27093,
         n27094, n27095, n27096, n27097, n27098, n27099, n27100, n27101,
         n27102, n27103, n27104, n27105, n27106, n27107, n27108, n27109,
         n27110, n27111, n27112, n27113, n27114, n27115, n27116, n27117,
         n27118, n27119, n27120, n27121, n27122, n27123, n27124, n27125,
         n27126, n27127, n27128, n27129, n27130, n27131, n27132, n27133,
         n27134, n27135, n27136, n27137, n27138, n27139, n27140, n27141,
         n27142, n27143, n27144, n27145, n27146, n27147, n27148, n27149,
         n27150, n27151, n27152, n27153, n27154, n27155, n27156, n27157,
         n27158, n27159, n27160, n27161, n27162, n27163, n27164, n27165,
         n27166, n27167, n27168, n27169, n27170, n27171, n27172, n27173,
         n27174, n27175, n27176, n27177, n27178, n27179, n27180, n27181,
         n27182, n27183, n27184, n27185, n27186, n27187, n27188, n27189,
         n27190, n27191, n27192, n27193, n27194, n27195, n27196, n27197,
         n27198, n27199, n27200, n27201, n27202, n27203, n27204, n27205,
         n27206, n27207, n27208, n27209, n27210, n27211, n27212, n27213,
         n27214, n27215, n27216, n27217, n27218, n27219, n27220, n27221,
         n27222, n27223, n27224, n27225, n27226, n27227, n27228, n27229,
         n27230, n27231, n27232, n27233, n27234, n27235, n27236, n27237,
         n27238, n27239, n27240, n27241, n27242, n27243, n27244, n27245,
         n27246, n27247, n27248, n27249, n27250, n27251, n27252, n27253,
         n27254, n27255, n27256, n27257, n27258, n27259, n27260, n27261,
         n27262, n27263, n27264, n27265, n27266, n27267, n27268, n27269,
         n27270, n27271, n27272, n27273, n27274, n27275, n27276, n27277,
         n27278, n27279, n27280, n27281, n27282, n27283, n27284, n27285,
         n27286, n27287, n27288, n27289, n27290, n27291, n27292, n27293,
         n27294, n27295, n27296, n27297, n27298, n27299, n27300, n27301,
         n27302, n27303, n27304, n27305, n27306, n27307, n27308, n27309,
         n27310, n27311, n27312, n27313, n27314, n27315, n27316, n27317,
         n27318, n27319, n27320, n27321, n27322, n27323, n27324, n27325,
         n27326, n27327, n27328, n27329, n27330, n27331, n27332, n27333,
         n27334, n27335, n27336, n27337, n27338, n27339, n27340, n27341,
         n27342, n27343, n27344, n27345, n27346, n27347, n27348, n27349,
         n27350, n27351, n27352, n27353, n27354, n27355, n27356, n27357,
         n27358, n27359, n27360, n27361, n27362, n27363, n27364, n27365,
         n27366, n27367, n27368, n27369, n27370, n27371, n27372, n27373,
         n27374, n27375, n27376, n27377, n27378, n27379, n27380, n27381,
         n27382, n27383, n27384, n27385, n27386, n27387, n27388, n27389,
         n27390, n27391, n27392, n27393, n27394, n27395, n27396, n27397,
         n27398, n27399, n27400, n27401, n27402, n27403, n27404, n27405,
         n27406, n27407, n27408, n27409, n27410, n27411, n27412, n27413,
         n27414, n27415, n27416, n27417, n27418, n27419, n27420, n27421,
         n27422, n27423, n27424, n27425, n27426, n27427, n27428, n27429,
         n27430, n27431, n27432, n27433, n27434, n27435, n27436, n27437,
         n27438, n27439, n27440, n27441, n27442, n27443, n27444, n27445,
         n27446, n27447, n27448, n27449, n27450, n27451, n27452, n27453,
         n27454, n27455, n27456, n27457, n27458, n27459, n27460, n27461,
         n27462, n27463, n27464, n27465, n27466, n27467, n27468, n27469,
         n27470, n27471, n27472, n27473, n27474, n27475, n27476, n27477,
         n27478, n27479, n27480, n27481, n27482, n27483, n27484, n27485,
         n27486, n27487, n27488, n27489, n27490, n27491, n27492, n27493,
         n27494, n27495, n27496, n27497, n27498, n27499, n27500, n27501,
         n27502, n27503, n27504, n27505, n27506, n27507, n27508, n27509,
         n27510, n27511, n27512, n27513, n27514, n27515, n27516, n27517,
         n27518, n27519, n27520, n27521, n27522, n27523, n27524, n27525,
         n27526, n27527, n27528, n27529, n27530, n27531, n27532, n27533,
         n27534, n27535, n27536, n27537, n27538, n27539, n27540, n27541,
         n27542, n27543, n27544, n27545, n27546, n27547, n27548, n27549,
         n27550, n27551, n27552, n27553, n27554, n27555, n27556, n27557,
         n27558, n27559, n27560, n27561, n27562, n27563, n27564, n27565,
         n27566, n27567, n27568, n27569, n27570, n27571, n27572, n27573,
         n27574, n27575, n27576, n27577, n27578, n27579, n27580, n27581,
         n27582, n27583, n27584, n27585, n27586, n27587, n27588, n27589,
         n27590, n27591, n27592, n27593, n27594, n27595, n27596, n27597,
         n27598, n27599, n27600, n27601, n27602, n27603, n27604, n27605,
         n27606, n27607, n27608, n27609, n27610, n27611, n27612, n27613,
         n27614, n27615, n27616, n27617, n27618, n27619, n27620, n27621,
         n27622, n27623, n27624, n27625, n27626, n27627, n27628, n27629,
         n27630, n27631, n27632, n27633, n27634, n27635, n27636, n27637,
         n27638, n27639, n27640, n27641, n27642, n27643, n27644, n27645,
         n27646, n27647, n27648, n27649, n27650, n27651, n27652, n27653,
         n27654, n27655, n27656, n27657, n27658, n27659, n27660, n27661,
         n27662, n27663, n27664, n27665, n27666, n27667, n27668, n27669,
         n27670, n27671, n27672, n27673, n27674, n27675, n27676, n27677,
         n27678, n27679, n27680, n27681, n27682, n27683, n27684, n27685,
         n27686, n27687, n27688, n27689, n27690, n27691, n27692, n27693,
         n27694, n27695, n27696, n27697, n27698, n27699, n27700, n27701,
         n27702, n27703, n27704, n27705, n27706, n27707, n27708, n27709,
         n27710, n27711, n27712, n27713, n27714, n27715, n27716, n27717,
         n27718, n27719, n27720, n27721, n27722, n27723, n27724, n27725,
         n27726, n27727, n27728, n27729, n27730, n27731, n27732, n27733,
         n27734, n27735, n27736, n27737, n27738, n27739, n27740, n27741,
         n27742, n27743, n27744, n27745, n27746, n27747, n27748, n27749,
         n27750, n27751, n27752, n27753, n27754, n27755, n27756, n27757,
         n27758, n27759, n27760, n27761, n27762, n27763, n27764, n27765,
         n27766, n27767, n27768, n27769, n27770, n27771, n27772, n27773,
         n27774, n27775, n27776, n27777, n27778, n27779, n27780, n27781,
         n27782, n27783, n27784, n27785, n27786, n27787, n27788, n27789,
         n27790, n27791, n27792, n27793, n27794, n27795, n27796, n27797,
         n27798, n27799, n27800, n27801, n27802, n27803, n27804, n27805,
         n27806, n27807, n27808, n27809, n27810, n27811, n27812, n27813,
         n27814, n27815, n27816, n27817, n27818, n27819, n27820, n27821,
         n27822, n27823, n27824, n27825, n27826, n27827, n27828, n27829,
         n27830, n27831, n27832, n27833, n27834, n27835, n27836, n27837,
         n27838, n27839, n27840, n27841, n27842, n27843, n27844, n27845,
         n27846, n27847, n27848, n27849, n27850, n27851, n27852, n27853,
         n27854, n27855, n27856, n27857, n27858, n27859, n27860, n27861,
         n27862, n27863, n27864, n27865, n27866, n27867, n27868, n27869,
         n27870, n27871, n27872, n27873, n27874, n27875, n27876, n27877,
         n27878, n27879, n27880, n27881, n27882, n27883, n27884, n27885,
         n27886, n27887, n27888, n27889, n27890, n27891, n27892, n27893,
         n27894, n27895, n27896, n27897, n27898, n27899, n27900, n27901,
         n27902, n27903, n27904, n27905, n27906, n27907, n27908, n27909,
         n27910, n27911, n27912, n27913, n27914, n27915, n27916, n27917,
         n27918, n27919, n27920, n27921, n27922, n27923, n27924, n27925,
         n27926, n27927, n27928, n27929, n27930, n27931, n27932, n27933,
         n27934, n27935, n27936, n27937, n27938, n27939, n27940, n27941,
         n27942, n27943, n27944, n27945, n27946, n27947, n27948, n27949,
         n27950, n27951, n27952, n27953, n27954, n27955, n27956, n27957,
         n27958, n27959, n27960, n27961, n27962, n27963, n27964, n27965,
         n27966, n27967, n27968, n27969, n27970, n27971, n27972, n27973,
         n27974, n27975, n27976, n27977, n27978, n27979, n27980, n27981,
         n27982, n27983, n27984, n27985, n27986, n27987, n27988, n27989,
         n27990, n27991, n27992, n27993, n27994, n27995, n27996, n27997,
         n27998, n27999, n28000, n28001, n28002, n28003, n28004, n28005,
         n28006, n28007, n28008, n28009, n28010, n28011, n28012, n28013,
         n28014, n28015, n28016, n28017, n28018, n28019, n28020, n28021,
         n28022, n28023, n28024, n28025, n28026, n28027, n28028, n28029,
         n28030, n28031, n28032, n28033, n28034, n28035, n28036, n28037,
         n28038, n28039, n28040, n28041, n28042, n28043, n28044, n28045,
         n28046, n28047, n28048, n28049, n28050, n28051, n28052, n28053,
         n28054, n28055, n28056, n28057, n28058, n28059, n28060, n28061,
         n28062, n28063, n28064, n28065, n28066, n28067, n28068, n28069,
         n28070, n28071, n28072, n28073, n28074, n28075, n28076, n28077,
         n28078, n28079, n28080, n28081, n28082, n28083, n28084, n28085,
         n28086, n28087, n28088, n28089, n28090, n28091, n28092, n28093,
         n28094, n28095, n28096, n28097, n28098, n28099, n28100, n28101,
         n28102, n28103, n28104, n28105, n28106, n28107, n28108, n28109,
         n28110, n28111, n28112, n28113, n28114, n28115, n28116, n28117,
         n28118, n28119, n28120, n28121, n28122, n28123, n28124, n28125,
         n28126, n28127, n28128, n28129, n28130, n28131, n28132, n28133,
         n28134, n28135, n28136, n28137, n28138, n28139, n28140, n28141,
         n28142, n28143, n28144, n28145, n28146, n28147, n28148, n28149,
         n28150, n28151, n28152, n28153, n28154, n28155, n28156, n28157,
         n28158, n28159, n28160, n28161, n28162, n28163, n28164, n28165,
         n28166, n28167, n28168, n28169, n28170, n28171, n28172, n28173,
         n28174, n28175, n28176, n28177, n28178, n28179, n28180, n28181,
         n28182, n28183, n28184, n28185, n28186, n28187, n28188, n28189,
         n28190, n28191, n28192, n28193, n28194, n28195, n28196, n28197,
         n28198, n28199, n28200, n28201, n28202, n28203, n28204, n28205,
         n28206, n28207, n28208, n28209, n28210, n28211, n28212, n28213,
         n28214, n28215, n28216, n28217, n28218, n28219, n28220, n28221,
         n28222, n28223, n28224, n28225, n28226, n28227, n28228, n28229,
         n28230, n28231, n28232, n28233, n28234, n28235, n28236, n28237,
         n28238, n28239, n28240, n28241, n28242, n28243, n28244, n28245,
         n28246, n28247, n28248, n28249, n28250, n28251, n28252, n28253,
         n28254, n28255, n28256, n28257, n28258, n28259, n28260, n28261,
         n28262, n28263, n28264, n28265, n28266, n28267, n28268, n28269,
         n28270, n28271, n28272, n28273, n28274, n28275, n28276, n28277,
         n28278, n28279, n28280, n28281, n28282, n28283, n28284, n28285,
         n28286, n28287, n28288, n28289, n28290, n28291, n28292, n28293,
         n28294, n28295, n28296, n28297, n28298, n28299, n28300, n28301,
         n28302, n28303, n28304, n28305, n28306, n28307, n28308, n28309,
         n28310, n28311, n28312, n28313, n28314, n28315, n28316, n28317,
         n28318, n28319, n28320, n28321, n28322, n28323, n28324, n28325,
         n28326, n28327, n28328, n28329, n28330, n28331, n28332, n28333,
         n28334, n28335, n28336, n28337, n28338, n28339, n28340, n28341,
         n28342, n28343, n28344, n28345, n28346, n28347, n28348, n28349,
         n28350, n28351, n28352, n28353, n28354, n28355, n28356, n28357,
         n28358, n28359, n28360, n28361, n28362, n28363, n28364, n28365,
         n28366, n28367, n28368, n28369, n28370, n28371, n28372, n28373,
         n28374, n28375, n28376, n28377, n28378, n28379, n28380, n28381,
         n28382, n28383, n28384, n28385, n28386, n28387, n28388, n28389,
         n28390, n28391, n28392, n28393, n28394, n28395, n28396, n28397,
         n28398, n28399, n28400, n28401, n28402, n28403, n28404, n28405,
         n28406, n28407, n28408, n28409, n28410, n28411, n28412, n28413,
         n28414, n28415, n28416, n28417, n28418, n28419, n28420, n28421,
         n28422, n28423, n28424, n28425, n28426, n28427, n28428, n28429,
         n28430, n28431, n28432, n28433, n28434, n28435, n28436, n28437,
         n28438, n28439, n28440, n28441, n28442, n28443, n28444, n28445,
         n28446, n28447, n28448, n28449, n28450, n28451, n28452, n28453,
         n28454, n28455, n28456, n28457, n28458, n28459, n28460, n28461,
         n28462, n28463, n28464, n28465, n28466, n28467, n28468, n28469,
         n28470, n28471, n28472, n28473, n28474, n28475, n28476, n28477,
         n28478, n28479, n28480, n28481, n28482, n28483, n28484, n28485,
         n28486, n28487, n28488, n28489, n28490, n28491, n28492, n28493,
         n28494, n28495, n28496, n28497, n28498, n28499, n28500, n28501,
         n28502, n28503, n28504, n28505, n28506, n28507, n28508, n28509,
         n28510, n28511, n28512, n28513, n28514, n28515, n28516, n28517,
         n28518, n28519, n28520, n28521, n28522, n28523, n28524, n28525,
         n28526, n28527, n28528, n28529, n28530, n28531, n28532, n28533,
         n28534, n28535, n28536, n28537, n28538, n28539, n28540, n28541,
         n28542, n28543, n28544, n28545, n28546, n28547, n28548, n28549,
         n28550, n28551, n28552, n28553, n28554, n28555, n28556, n28557,
         n28558, n28559, n28560, n28561, n28562, n28563, n28564, n28565,
         n28566, n28567, n28568, n28569, n28570, n28571, n28572, n28573,
         n28574, n28575, n28576, n28577, n28578, n28579, n28580, n28581,
         n28582, n28583, n28584, n28585, n28586, n28587, n28588, n28589,
         n28590, n28591, n28592, n28593, n28594, n28595, n28596, n28597,
         n28598, n28599, n28600, n28601, n28602, n28603, n28604, n28605,
         n28606, n28607, n28608, n28609, n28610, n28611, n28612, n28613,
         n28614, n28615, n28616, n28617, n28618, n28619, n28620, n28621,
         n28622, n28623, n28624, n28625, n28626, n28627, n28628, n28629,
         n28630, n28631, n28632, n28633, n28634, n28635, n28636, n28637,
         n28638, n28639, n28640, n28641, n28642, n28643, n28644, n28645,
         n28646, n28647, n28648, n28649, n28650, n28651, n28652, n28653,
         n28654, n28655, n28656, n28657, n28658, n28659, n28660, n28661,
         n28662, n28663, n28664, n28665, n28666, n28667, n28668, n28669,
         n28670, n28671, n28672, n28673, n28674, n28675, n28676, n28677,
         n28678, n28679, n28680, n28681, n28682, n28683, n28684, n28685,
         n28686, n28687, n28688, n28689, n28690, n28691, n28692, n28693,
         n28694, n28695, n28696, n28697, n28698, n28699, n28700, n28701,
         n28702, n28703, n28704, n28705, n28706, n28707, n28708, n28709,
         n28710, n28711, n28712, n28713, n28714, n28715, n28716, n28717,
         n28718, n28719, n28720, n28721, n28722, n28723, n28724, n28725,
         n28726, n28727, n28728, n28729, n28730, n28731, n28732, n28733,
         n28734, n28735, n28736, n28737, n28738, n28739, n28740, n28741,
         n28742, n28743, n28744, n28745, n28746, n28747, n28748, n28749,
         n28750, n28751, n28752, n28753, n28754, n28755, n28756, n28757,
         n28758, n28759, n28760, n28761, n28762, n28763, n28764, n28765,
         n28766, n28767, n28768, n28769, n28770, n28771, n28772, n28773,
         n28774, n28775, n28776, n28777, n28778, n28779, n28780, n28781,
         n28782, n28783, n28784, n28785, n28786, n28787, n28788, n28789,
         n28790, n28791, n28792, n28793, n28794, n28795, n28796, n28797,
         n28798, n28799, n28800, n28801, n28802, n28803, n28804, n28805,
         n28806, n28807, n28808, n28809, n28810, n28811, n28812, n28813,
         n28814, n28815, n28816, n28817, n28818, n28819, n28820, n28821,
         n28822, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5;
  wire   [618:604] n;
  wire   [5:2] add_283_carry;
  wire   [9:2] add_262_carry;
  assign dut__dim__address[8] = 1'b0;
  assign dut__dim__write = 1'b0;
  assign dut__bvm__write = 1'b0;
  assign dut__dim__enable = 1'b1;

  macopertion_1 W ( .in_a_mac({n4967, n4966, n4965, n4964, n4963, n4962, n4961, 
        n4960, n4959, n4958, n4957, n4956, n4955, n4954, n4953, n4952}), 
        .in_b_mac({n25960, n25962, n25964, n25966, n25968, n25970, n25972, 
        n25974, n25975, n25977, n25978, n25979, n25769, n25981, n25754, n4888}), .bitselect1({add_180_A_3_, add_180_A_2_, add_180_A_1_, add_180_A_0_}), .clk(
        clk), .min({SYNOPSYS_UNCONNECTED_1, n2401, n2400, n2399, n2398, n2397, 
        n2396, n2395, n2394, n2393, n2392, n2391, n2390, n2389, n2388, n2387})
         );
  macopertion_3 X ( .in_a_mac({n4951, n4950, n4949, n4948, n4947, n4946, n4945, 
        n4944, n4943, n4942, n4941, n4940, n4939, n4938, n4937, n4936}), 
        .in_b_mac({n25960, n25962, n25964, n25966, n25968, n25970, n25972, 
        n25974, n25975, n25977, n25978, n25979, n25769, n25981, n25754, n4888}), .bitselect1({add_180_A_3_, add_180_A_2_, add_180_A_1_, add_180_A_0_}), .clk(
        clk), .min({SYNOPSYS_UNCONNECTED_2, n2385, n2384, n2383, n2382, n2381, 
        n2380, n2379, n2378, n2377, n2376, n2375, n2374, n2373, n2372, n2371})
         );
  macopertion_2 Y ( .in_a_mac({n4935, n4934, n4933, n4932, n4931, n4930, n4929, 
        n4928, n4927, n4926, n4925, n4924, n4923, n4922, n4921, n4920}), 
        .in_b_mac({n25960, n25962, n25964, n25966, n25968, n25970, n25972, 
        n25974, n25975, n25977, n25978, n25979, n25732, n25981, n25754, n4888}), .bitselect1({add_180_A_3_, add_180_A_2_, add_180_A_1_, add_180_A_0_}), .clk(
        clk), .min({SYNOPSYS_UNCONNECTED_3, n2369, n2368, n2367, n2366, n2365, 
        n2364, n2363, n2362, n2361, n2360, n2359, n2358, n2357, n2356, n2355})
         );
  macopertion_0 Z ( .in_a_mac({n4919, n4918, n4917, n4916, n4915, n4914, n4913, 
        n4912, n25751, n4910, n25780, n25762, n25765, n4906, n25763, n25752}), 
        .in_b_mac({n25960, n25962, n25964, n25966, n25968, n25970, n25972, 
        n25974, n25975, n25977, n25978, n25741, n25980, n25761, n25983, n4888}), .bitselect1({add_180_A_3_, add_180_A_2_, add_180_A_1_, add_180_A_0_}), .clk(
        clk), .min({SYNOPSYS_UNCONNECTED_4, n2353, n2352, n2351, n2350, n2349, 
        n2348, n2347, n2346, n2345, n2344, n2343, n2342, n2341, n2340, n2339})
         );
  macopertion_m Z1 ( .in_z_mac({n651, n650, n649, n648, n647, n646, n645, n644, 
        n643, n642, n25766, n25759, n25764, n25747, n25767, n636}), .in_m_mac(
        {n5056, n5055, n5054, n5053, n5052, n5051, n5050, n5049, n5048, n5047, 
        n25738, n25748, n25779, n25737, n25760, n5041}), .sendz_count({
        add_283_A_5_, add_283_A_4_, add_283_A_3_, add_283_A_2_, add_283_A_1_, 
        add_283_A_0_}), .clk(clk), .minm({SYNOPSYS_UNCONNECTED_5, n}) );
  HA_X1 add_262_U1_1_1 ( .A(add_1445_B_1_), .B(add_1445_B_0_), .CO(
        add_262_carry[2]), .S(U8_DATA2_1) );
  HA_X1 add_262_U1_1_2 ( .A(add_1445_B_2_), .B(add_262_carry[2]), .CO(
        add_262_carry[3]), .S(U8_DATA2_2) );
  HA_X1 add_262_U1_1_3 ( .A(add_1445_B_3_), .B(add_262_carry[3]), .CO(
        add_262_carry[4]), .S(U8_DATA2_3) );
  HA_X1 add_262_U1_1_4 ( .A(add_1445_B_4_), .B(add_262_carry[4]), .CO(
        add_262_carry[5]), .S(U8_DATA2_4) );
  HA_X1 add_262_U1_1_5 ( .A(add_1445_B_5_), .B(add_262_carry[5]), .CO(
        add_262_carry[6]), .S(U8_DATA2_5) );
  HA_X1 add_262_U1_1_6 ( .A(add_1445_B_6_), .B(add_262_carry[6]), .CO(
        add_262_carry[7]), .S(U8_DATA2_6) );
  HA_X1 add_262_U1_1_7 ( .A(add_1445_B_7_), .B(add_262_carry[7]), .CO(
        add_262_carry[8]), .S(U8_DATA2_7) );
  HA_X1 add_262_U1_1_8 ( .A(add_1445_B_8_), .B(add_262_carry[8]), .CO(
        add_262_carry[9]), .S(U8_DATA2_8) );
  HA_X1 add_283_U1_1_1 ( .A(add_283_A_1_), .B(add_283_A_0_), .CO(
        add_283_carry[2]), .S(U7_DATA2_1) );
  HA_X1 add_283_U1_1_2 ( .A(add_283_A_2_), .B(add_283_carry[2]), .CO(
        add_283_carry[3]), .S(U7_DATA2_2) );
  HA_X1 add_283_U1_1_3 ( .A(add_283_A_3_), .B(add_283_carry[3]), .CO(
        add_283_carry[4]), .S(U7_DATA2_3) );
  HA_X1 add_283_U1_1_4 ( .A(add_283_A_4_), .B(add_283_carry[4]), .CO(
        add_283_carry[5]), .S(U7_DATA2_4) );
  DFF_X1 flag_out_reg ( .D(n24823), .CK(clk), .QN(n22427) );
  DFF_X1 count_store_reg_1_ ( .D(n24821), .CK(clk), .Q(n24891), .QN(n22423) );
  DFF_X1 count_store_reg_2_ ( .D(n24820), .CK(clk), .Q(n25248), .QN(n22422) );
  DFF_X1 count_store_reg_0_ ( .D(n24822), .CK(clk), .Q(n24868), .QN(n22424) );
  DFF_X1 bitselect_reg_0_ ( .D(n24817), .CK(clk), .Q(n24833), .QN(n22386) );
  DFF_X1 bitselect_reg_1_ ( .D(n24816), .CK(clk), .Q(n25400), .QN(n22385) );
  DFF_X1 counter_reg_0_ ( .D(n24813), .CK(clk), .Q(n25254), .QN(n22390) );
  DFF_X1 counter_reg_1_ ( .D(n24812), .CK(clk), .Q(n25256), .QN(n22389) );
  DFF_X1 counter_reg_2_ ( .D(n24811), .CK(clk), .Q(n25252), .QN(n22388) );
  DFF_X1 counter_reg_3_ ( .D(n24810), .CK(clk), .Q(n24895), .QN(n22387) );
  DFF_X1 bitselect_reg_2_ ( .D(n24815), .CK(clk), .Q(n24832), .QN(n22384) );
  DFF_X1 bitselect_reg_3_ ( .D(n24814), .CK(clk), .Q(n25249), .QN(n22383) );
  DFF_X1 avector23_reg_5__0_ ( .D(n22380), .CK(clk), .QN(n17557) );
  DFF_X1 avector23_reg_5__1_ ( .D(n22379), .CK(clk), .QN(n17520) );
  DFF_X1 avector23_reg_5__2_ ( .D(n22378), .CK(clk), .QN(n17483) );
  DFF_X1 avector23_reg_5__3_ ( .D(n22377), .CK(clk), .QN(n17446) );
  DFF_X1 avector23_reg_5__4_ ( .D(n22376), .CK(clk), .QN(n17409) );
  DFF_X1 avector23_reg_5__5_ ( .D(n22375), .CK(clk), .QN(n17372) );
  DFF_X1 avector23_reg_5__6_ ( .D(n22374), .CK(clk), .QN(n17335) );
  DFF_X1 avector23_reg_5__7_ ( .D(n22373), .CK(clk), .QN(n17298) );
  DFF_X1 avector23_reg_5__8_ ( .D(n22372), .CK(clk), .QN(n17261) );
  DFF_X1 avector23_reg_5__9_ ( .D(n22371), .CK(clk), .QN(n17224) );
  DFF_X1 avector23_reg_5__10_ ( .D(n22370), .CK(clk), .QN(n17187) );
  DFF_X1 avector23_reg_5__11_ ( .D(n22369), .CK(clk), .QN(n17150) );
  DFF_X1 avector23_reg_5__12_ ( .D(n22368), .CK(clk), .QN(n17113) );
  DFF_X1 avector23_reg_5__13_ ( .D(n22367), .CK(clk), .QN(n17076) );
  DFF_X1 avector23_reg_5__14_ ( .D(n22366), .CK(clk), .QN(n17039) );
  DFF_X1 avector23_reg_5__15_ ( .D(n22365), .CK(clk), .QN(n17002) );
  DFF_X1 avector13_reg_5__0_ ( .D(n22316), .CK(clk), .QN(n18149) );
  DFF_X1 avector13_reg_5__1_ ( .D(n22315), .CK(clk), .QN(n18112) );
  DFF_X1 avector13_reg_5__2_ ( .D(n22314), .CK(clk), .QN(n18075) );
  DFF_X1 avector13_reg_5__3_ ( .D(n22313), .CK(clk), .QN(n18038) );
  DFF_X1 avector13_reg_5__4_ ( .D(n22312), .CK(clk), .QN(n18001) );
  DFF_X1 avector13_reg_5__5_ ( .D(n22311), .CK(clk), .QN(n17964) );
  DFF_X1 avector13_reg_5__6_ ( .D(n22310), .CK(clk), .QN(n17927) );
  DFF_X1 avector13_reg_5__7_ ( .D(n22309), .CK(clk), .QN(n17890) );
  DFF_X1 avector13_reg_5__8_ ( .D(n22308), .CK(clk), .QN(n17853) );
  DFF_X1 avector13_reg_5__9_ ( .D(n22307), .CK(clk), .QN(n17816) );
  DFF_X1 avector13_reg_5__10_ ( .D(n22306), .CK(clk), .QN(n17779) );
  DFF_X1 avector13_reg_5__11_ ( .D(n22305), .CK(clk), .QN(n17742) );
  DFF_X1 avector13_reg_5__12_ ( .D(n22304), .CK(clk), .QN(n17705) );
  DFF_X1 avector13_reg_5__13_ ( .D(n22303), .CK(clk), .QN(n17668) );
  DFF_X1 avector13_reg_5__14_ ( .D(n22302), .CK(clk), .QN(n17631) );
  DFF_X1 avector13_reg_5__15_ ( .D(n22301), .CK(clk), .QN(n17594) );
  DFF_X1 avector03_reg_5__0_ ( .D(n22252), .CK(clk), .QN(n18741) );
  DFF_X1 avector03_reg_5__1_ ( .D(n22251), .CK(clk), .QN(n18704) );
  DFF_X1 avector03_reg_5__2_ ( .D(n22250), .CK(clk), .QN(n18667) );
  DFF_X1 avector03_reg_5__3_ ( .D(n22249), .CK(clk), .QN(n18630) );
  DFF_X1 avector03_reg_5__4_ ( .D(n22248), .CK(clk), .QN(n18593) );
  DFF_X1 avector03_reg_5__5_ ( .D(n22247), .CK(clk), .QN(n18556) );
  DFF_X1 avector03_reg_5__6_ ( .D(n22246), .CK(clk), .QN(n18519) );
  DFF_X1 avector03_reg_5__7_ ( .D(n22245), .CK(clk), .QN(n18482) );
  DFF_X1 avector03_reg_5__8_ ( .D(n22244), .CK(clk), .QN(n18445) );
  DFF_X1 avector03_reg_5__9_ ( .D(n22243), .CK(clk), .QN(n18408) );
  DFF_X1 avector03_reg_5__10_ ( .D(n22242), .CK(clk), .QN(n18371) );
  DFF_X1 avector03_reg_5__11_ ( .D(n22241), .CK(clk), .QN(n18334) );
  DFF_X1 avector03_reg_5__12_ ( .D(n22240), .CK(clk), .QN(n18297) );
  DFF_X1 avector03_reg_5__13_ ( .D(n22239), .CK(clk), .QN(n18260) );
  DFF_X1 avector03_reg_5__14_ ( .D(n22238), .CK(clk), .QN(n18223) );
  DFF_X1 avector03_reg_5__15_ ( .D(n22237), .CK(clk), .QN(n18186) );
  DFF_X1 avector33_reg_5__0_ ( .D(n21148), .CK(clk), .QN(n16965) );
  DFF_X1 avector33_reg_5__1_ ( .D(n21147), .CK(clk), .QN(n16928) );
  DFF_X1 avector33_reg_5__2_ ( .D(n21146), .CK(clk), .QN(n16891) );
  DFF_X1 avector33_reg_5__3_ ( .D(n21145), .CK(clk), .QN(n16854) );
  DFF_X1 avector33_reg_5__4_ ( .D(n21144), .CK(clk), .QN(n16817) );
  DFF_X1 avector33_reg_5__5_ ( .D(n21143), .CK(clk), .QN(n16780) );
  DFF_X1 avector33_reg_5__6_ ( .D(n21142), .CK(clk), .QN(n16743) );
  DFF_X1 avector33_reg_5__7_ ( .D(n21141), .CK(clk), .QN(n16706) );
  DFF_X1 avector33_reg_5__8_ ( .D(n21140), .CK(clk), .QN(n16669) );
  DFF_X1 avector33_reg_5__9_ ( .D(n21139), .CK(clk), .QN(n16632) );
  DFF_X1 avector33_reg_5__10_ ( .D(n21138), .CK(clk), .QN(n16595) );
  DFF_X1 avector33_reg_5__11_ ( .D(n21137), .CK(clk), .QN(n16558) );
  DFF_X1 avector33_reg_5__12_ ( .D(n21136), .CK(clk), .QN(n16521) );
  DFF_X1 avector33_reg_5__13_ ( .D(n21135), .CK(clk), .QN(n16484) );
  DFF_X1 avector33_reg_5__14_ ( .D(n21134), .CK(clk), .QN(n16447) );
  DFF_X1 avector33_reg_5__15_ ( .D(n21133), .CK(clk), .QN(n16410) );
  DFF_X1 avector22_reg_5__0_ ( .D(n22188), .CK(clk), .QN(n17530) );
  DFF_X1 avector22_reg_5__1_ ( .D(n22187), .CK(clk), .QN(n17493) );
  DFF_X1 avector22_reg_5__2_ ( .D(n22186), .CK(clk), .QN(n17456) );
  DFF_X1 avector22_reg_5__3_ ( .D(n22185), .CK(clk), .QN(n17419) );
  DFF_X1 avector22_reg_5__4_ ( .D(n22184), .CK(clk), .QN(n17382) );
  DFF_X1 avector22_reg_5__5_ ( .D(n22183), .CK(clk), .QN(n17345) );
  DFF_X1 avector22_reg_5__6_ ( .D(n22182), .CK(clk), .QN(n17308) );
  DFF_X1 avector22_reg_5__7_ ( .D(n22181), .CK(clk), .QN(n17271) );
  DFF_X1 avector22_reg_5__8_ ( .D(n22180), .CK(clk), .QN(n17234) );
  DFF_X1 avector22_reg_5__9_ ( .D(n22179), .CK(clk), .QN(n17197) );
  DFF_X1 avector22_reg_5__10_ ( .D(n22178), .CK(clk), .QN(n17160) );
  DFF_X1 avector22_reg_5__11_ ( .D(n22177), .CK(clk), .QN(n17123) );
  DFF_X1 avector22_reg_5__12_ ( .D(n22176), .CK(clk), .QN(n17086) );
  DFF_X1 avector22_reg_5__13_ ( .D(n22175), .CK(clk), .QN(n17049) );
  DFF_X1 avector22_reg_5__14_ ( .D(n22174), .CK(clk), .QN(n17012) );
  DFF_X1 avector22_reg_5__15_ ( .D(n22173), .CK(clk), .QN(n16975) );
  DFF_X1 avector12_reg_5__0_ ( .D(n22124), .CK(clk), .QN(n18122) );
  DFF_X1 avector12_reg_5__1_ ( .D(n22123), .CK(clk), .QN(n18085) );
  DFF_X1 avector12_reg_5__2_ ( .D(n22122), .CK(clk), .QN(n18048) );
  DFF_X1 avector12_reg_5__3_ ( .D(n22121), .CK(clk), .QN(n18011) );
  DFF_X1 avector12_reg_5__4_ ( .D(n22120), .CK(clk), .QN(n17974) );
  DFF_X1 avector12_reg_5__5_ ( .D(n22119), .CK(clk), .QN(n17937) );
  DFF_X1 avector12_reg_5__6_ ( .D(n22118), .CK(clk), .QN(n17900) );
  DFF_X1 avector12_reg_5__7_ ( .D(n22117), .CK(clk), .QN(n17863) );
  DFF_X1 avector12_reg_5__8_ ( .D(n22116), .CK(clk), .QN(n17826) );
  DFF_X1 avector12_reg_5__9_ ( .D(n22115), .CK(clk), .QN(n17789) );
  DFF_X1 avector12_reg_5__10_ ( .D(n22114), .CK(clk), .QN(n17752) );
  DFF_X1 avector12_reg_5__11_ ( .D(n22113), .CK(clk), .QN(n17715) );
  DFF_X1 avector12_reg_5__12_ ( .D(n22112), .CK(clk), .QN(n17678) );
  DFF_X1 avector12_reg_5__13_ ( .D(n22111), .CK(clk), .QN(n17641) );
  DFF_X1 avector12_reg_5__14_ ( .D(n22110), .CK(clk), .QN(n17604) );
  DFF_X1 avector12_reg_5__15_ ( .D(n22109), .CK(clk), .QN(n17567) );
  DFF_X1 avector02_reg_5__0_ ( .D(n22060), .CK(clk), .QN(n18714) );
  DFF_X1 avector02_reg_5__1_ ( .D(n22059), .CK(clk), .QN(n18677) );
  DFF_X1 avector02_reg_5__2_ ( .D(n22058), .CK(clk), .QN(n18640) );
  DFF_X1 avector02_reg_5__3_ ( .D(n22057), .CK(clk), .QN(n18603) );
  DFF_X1 avector02_reg_5__4_ ( .D(n22056), .CK(clk), .QN(n18566) );
  DFF_X1 avector02_reg_5__5_ ( .D(n22055), .CK(clk), .QN(n18529) );
  DFF_X1 avector02_reg_5__6_ ( .D(n22054), .CK(clk), .QN(n18492) );
  DFF_X1 avector02_reg_5__7_ ( .D(n22053), .CK(clk), .QN(n18455) );
  DFF_X1 avector02_reg_5__8_ ( .D(n22052), .CK(clk), .QN(n18418) );
  DFF_X1 avector02_reg_5__9_ ( .D(n22051), .CK(clk), .QN(n18381) );
  DFF_X1 avector02_reg_5__10_ ( .D(n22050), .CK(clk), .QN(n18344) );
  DFF_X1 avector02_reg_5__11_ ( .D(n22049), .CK(clk), .QN(n18307) );
  DFF_X1 avector02_reg_5__12_ ( .D(n22048), .CK(clk), .QN(n18270) );
  DFF_X1 avector02_reg_5__13_ ( .D(n22047), .CK(clk), .QN(n18233) );
  DFF_X1 avector02_reg_5__14_ ( .D(n22046), .CK(clk), .QN(n18196) );
  DFF_X1 avector02_reg_5__15_ ( .D(n22045), .CK(clk), .QN(n18159) );
  DFF_X1 avector32_reg_5__0_ ( .D(n21996), .CK(clk), .QN(n16938) );
  DFF_X1 avector32_reg_5__1_ ( .D(n21995), .CK(clk), .QN(n16901) );
  DFF_X1 avector32_reg_5__2_ ( .D(n21994), .CK(clk), .QN(n16864) );
  DFF_X1 avector32_reg_5__3_ ( .D(n21993), .CK(clk), .QN(n16827) );
  DFF_X1 avector32_reg_5__4_ ( .D(n21992), .CK(clk), .QN(n16790) );
  DFF_X1 avector32_reg_5__5_ ( .D(n21991), .CK(clk), .QN(n16753) );
  DFF_X1 avector32_reg_5__6_ ( .D(n21990), .CK(clk), .QN(n16716) );
  DFF_X1 avector32_reg_5__7_ ( .D(n21989), .CK(clk), .QN(n16679) );
  DFF_X1 avector32_reg_5__8_ ( .D(n21988), .CK(clk), .QN(n16642) );
  DFF_X1 avector32_reg_5__9_ ( .D(n21987), .CK(clk), .QN(n16605) );
  DFF_X1 avector32_reg_5__10_ ( .D(n21986), .CK(clk), .QN(n16568) );
  DFF_X1 avector32_reg_5__11_ ( .D(n21985), .CK(clk), .QN(n16531) );
  DFF_X1 avector32_reg_5__12_ ( .D(n21984), .CK(clk), .QN(n16494) );
  DFF_X1 avector32_reg_5__13_ ( .D(n21983), .CK(clk), .QN(n16457) );
  DFF_X1 avector32_reg_5__14_ ( .D(n21982), .CK(clk), .QN(n16420) );
  DFF_X1 avector32_reg_5__15_ ( .D(n21981), .CK(clk), .QN(n16383) );
  DFF_X1 avector21_reg_5__0_ ( .D(n21932), .CK(clk), .QN(n17539) );
  DFF_X1 avector21_reg_5__1_ ( .D(n21931), .CK(clk), .QN(n17502) );
  DFF_X1 avector21_reg_5__2_ ( .D(n21930), .CK(clk), .QN(n17465) );
  DFF_X1 avector21_reg_5__3_ ( .D(n21929), .CK(clk), .QN(n17428) );
  DFF_X1 avector21_reg_5__4_ ( .D(n21928), .CK(clk), .QN(n17391) );
  DFF_X1 avector21_reg_5__5_ ( .D(n21927), .CK(clk), .QN(n17354) );
  DFF_X1 avector21_reg_5__6_ ( .D(n21926), .CK(clk), .QN(n17317) );
  DFF_X1 avector21_reg_5__7_ ( .D(n21925), .CK(clk), .QN(n17280) );
  DFF_X1 avector21_reg_5__8_ ( .D(n21924), .CK(clk), .QN(n17243) );
  DFF_X1 avector21_reg_5__9_ ( .D(n21923), .CK(clk), .QN(n17206) );
  DFF_X1 avector21_reg_5__10_ ( .D(n21922), .CK(clk), .QN(n17169) );
  DFF_X1 avector21_reg_5__11_ ( .D(n21921), .CK(clk), .QN(n17132) );
  DFF_X1 avector21_reg_5__12_ ( .D(n21920), .CK(clk), .QN(n17095) );
  DFF_X1 avector21_reg_5__13_ ( .D(n21919), .CK(clk), .QN(n17058) );
  DFF_X1 avector21_reg_5__14_ ( .D(n21918), .CK(clk), .QN(n17021) );
  DFF_X1 avector21_reg_5__15_ ( .D(n21917), .CK(clk), .QN(n16984) );
  DFF_X1 avector11_reg_5__0_ ( .D(n21868), .CK(clk), .QN(n18131) );
  DFF_X1 avector11_reg_5__1_ ( .D(n21867), .CK(clk), .QN(n18094) );
  DFF_X1 avector11_reg_5__2_ ( .D(n21866), .CK(clk), .QN(n18057) );
  DFF_X1 avector11_reg_5__3_ ( .D(n21865), .CK(clk), .QN(n18020) );
  DFF_X1 avector11_reg_5__4_ ( .D(n21864), .CK(clk), .QN(n17983) );
  DFF_X1 avector11_reg_5__5_ ( .D(n21863), .CK(clk), .QN(n17946) );
  DFF_X1 avector11_reg_5__6_ ( .D(n21862), .CK(clk), .QN(n17909) );
  DFF_X1 avector11_reg_5__7_ ( .D(n21861), .CK(clk), .QN(n17872) );
  DFF_X1 avector11_reg_5__8_ ( .D(n21860), .CK(clk), .QN(n17835) );
  DFF_X1 avector11_reg_5__9_ ( .D(n21859), .CK(clk), .QN(n17798) );
  DFF_X1 avector11_reg_5__10_ ( .D(n21858), .CK(clk), .QN(n17761) );
  DFF_X1 avector11_reg_5__11_ ( .D(n21857), .CK(clk), .QN(n17724) );
  DFF_X1 avector11_reg_5__12_ ( .D(n21856), .CK(clk), .QN(n17687) );
  DFF_X1 avector11_reg_5__13_ ( .D(n21855), .CK(clk), .QN(n17650) );
  DFF_X1 avector11_reg_5__14_ ( .D(n21854), .CK(clk), .QN(n17613) );
  DFF_X1 avector11_reg_5__15_ ( .D(n21853), .CK(clk), .QN(n17576) );
  DFF_X1 avector01_reg_5__0_ ( .D(n21804), .CK(clk), .QN(n18723) );
  DFF_X1 avector01_reg_5__1_ ( .D(n21803), .CK(clk), .QN(n18686) );
  DFF_X1 avector01_reg_5__2_ ( .D(n21802), .CK(clk), .QN(n18649) );
  DFF_X1 avector01_reg_5__3_ ( .D(n21801), .CK(clk), .QN(n18612) );
  DFF_X1 avector01_reg_5__4_ ( .D(n21800), .CK(clk), .QN(n18575) );
  DFF_X1 avector01_reg_5__5_ ( .D(n21799), .CK(clk), .QN(n18538) );
  DFF_X1 avector01_reg_5__6_ ( .D(n21798), .CK(clk), .QN(n18501) );
  DFF_X1 avector01_reg_5__7_ ( .D(n21797), .CK(clk), .QN(n18464) );
  DFF_X1 avector01_reg_5__8_ ( .D(n21796), .CK(clk), .QN(n18427) );
  DFF_X1 avector01_reg_5__9_ ( .D(n21795), .CK(clk), .QN(n18390) );
  DFF_X1 avector01_reg_5__10_ ( .D(n21794), .CK(clk), .QN(n18353) );
  DFF_X1 avector01_reg_5__11_ ( .D(n21793), .CK(clk), .QN(n18316) );
  DFF_X1 avector01_reg_5__12_ ( .D(n21792), .CK(clk), .QN(n18279) );
  DFF_X1 avector01_reg_5__13_ ( .D(n21791), .CK(clk), .QN(n18242) );
  DFF_X1 avector01_reg_5__14_ ( .D(n21790), .CK(clk), .QN(n18205) );
  DFF_X1 avector01_reg_5__15_ ( .D(n21789), .CK(clk), .QN(n18168) );
  DFF_X1 avector31_reg_5__0_ ( .D(n21740), .CK(clk), .QN(n16947) );
  DFF_X1 avector31_reg_5__1_ ( .D(n21739), .CK(clk), .QN(n16910) );
  DFF_X1 avector31_reg_5__2_ ( .D(n21738), .CK(clk), .QN(n16873) );
  DFF_X1 avector31_reg_5__3_ ( .D(n21737), .CK(clk), .QN(n16836) );
  DFF_X1 avector31_reg_5__4_ ( .D(n21736), .CK(clk), .QN(n16799) );
  DFF_X1 avector31_reg_5__5_ ( .D(n21735), .CK(clk), .QN(n16762) );
  DFF_X1 avector31_reg_5__6_ ( .D(n21734), .CK(clk), .QN(n16725) );
  DFF_X1 avector31_reg_5__7_ ( .D(n21733), .CK(clk), .QN(n16688) );
  DFF_X1 avector31_reg_5__8_ ( .D(n21732), .CK(clk), .QN(n16651) );
  DFF_X1 avector31_reg_5__9_ ( .D(n21731), .CK(clk), .QN(n16614) );
  DFF_X1 avector31_reg_5__10_ ( .D(n21730), .CK(clk), .QN(n16577) );
  DFF_X1 avector31_reg_5__11_ ( .D(n21729), .CK(clk), .QN(n16540) );
  DFF_X1 avector31_reg_5__12_ ( .D(n21728), .CK(clk), .QN(n16503) );
  DFF_X1 avector31_reg_5__13_ ( .D(n21727), .CK(clk), .QN(n16466) );
  DFF_X1 avector31_reg_5__14_ ( .D(n21726), .CK(clk), .QN(n16429) );
  DFF_X1 avector31_reg_5__15_ ( .D(n21725), .CK(clk), .QN(n16392) );
  DFF_X1 avector20_reg_5__0_ ( .D(n21676), .CK(clk), .QN(n17548) );
  DFF_X1 avector20_reg_5__1_ ( .D(n21675), .CK(clk), .QN(n17511) );
  DFF_X1 avector20_reg_5__2_ ( .D(n21674), .CK(clk), .QN(n17474) );
  DFF_X1 avector20_reg_5__3_ ( .D(n21673), .CK(clk), .QN(n17437) );
  DFF_X1 avector20_reg_5__4_ ( .D(n21672), .CK(clk), .QN(n17400) );
  DFF_X1 avector20_reg_5__5_ ( .D(n21671), .CK(clk), .QN(n17363) );
  DFF_X1 avector20_reg_5__6_ ( .D(n21670), .CK(clk), .QN(n17326) );
  DFF_X1 avector20_reg_5__7_ ( .D(n21669), .CK(clk), .QN(n17289) );
  DFF_X1 avector20_reg_5__8_ ( .D(n21668), .CK(clk), .QN(n17252) );
  DFF_X1 avector20_reg_5__9_ ( .D(n21667), .CK(clk), .QN(n17215) );
  DFF_X1 avector20_reg_5__10_ ( .D(n21666), .CK(clk), .QN(n17178) );
  DFF_X1 avector20_reg_5__11_ ( .D(n21665), .CK(clk), .QN(n17141) );
  DFF_X1 avector20_reg_5__12_ ( .D(n21664), .CK(clk), .QN(n17104) );
  DFF_X1 avector20_reg_5__13_ ( .D(n21663), .CK(clk), .QN(n17067) );
  DFF_X1 avector20_reg_5__14_ ( .D(n21662), .CK(clk), .QN(n17030) );
  DFF_X1 avector20_reg_5__15_ ( .D(n21661), .CK(clk), .QN(n16993) );
  DFF_X1 avector10_reg_5__0_ ( .D(n21612), .CK(clk), .QN(n18140) );
  DFF_X1 avector10_reg_5__1_ ( .D(n21611), .CK(clk), .QN(n18103) );
  DFF_X1 avector10_reg_5__2_ ( .D(n21610), .CK(clk), .QN(n18066) );
  DFF_X1 avector10_reg_5__3_ ( .D(n21609), .CK(clk), .QN(n18029) );
  DFF_X1 avector10_reg_5__4_ ( .D(n21608), .CK(clk), .QN(n17992) );
  DFF_X1 avector10_reg_5__5_ ( .D(n21607), .CK(clk), .QN(n17955) );
  DFF_X1 avector10_reg_5__6_ ( .D(n21606), .CK(clk), .QN(n17918) );
  DFF_X1 avector10_reg_5__7_ ( .D(n21605), .CK(clk), .QN(n17881) );
  DFF_X1 avector10_reg_5__8_ ( .D(n21604), .CK(clk), .QN(n17844) );
  DFF_X1 avector10_reg_5__9_ ( .D(n21603), .CK(clk), .QN(n17807) );
  DFF_X1 avector10_reg_5__10_ ( .D(n21602), .CK(clk), .QN(n17770) );
  DFF_X1 avector10_reg_5__11_ ( .D(n21601), .CK(clk), .QN(n17733) );
  DFF_X1 avector10_reg_5__12_ ( .D(n21600), .CK(clk), .QN(n17696) );
  DFF_X1 avector10_reg_5__13_ ( .D(n21599), .CK(clk), .QN(n17659) );
  DFF_X1 avector10_reg_5__14_ ( .D(n21598), .CK(clk), .QN(n17622) );
  DFF_X1 avector10_reg_5__15_ ( .D(n21597), .CK(clk), .QN(n17585) );
  DFF_X1 avector00_reg_5__0_ ( .D(n21548), .CK(clk), .QN(n18732) );
  DFF_X1 avector00_reg_5__1_ ( .D(n21547), .CK(clk), .QN(n18695) );
  DFF_X1 avector00_reg_5__2_ ( .D(n21546), .CK(clk), .QN(n18658) );
  DFF_X1 avector00_reg_5__3_ ( .D(n21545), .CK(clk), .QN(n18621) );
  DFF_X1 avector00_reg_5__4_ ( .D(n21544), .CK(clk), .QN(n18584) );
  DFF_X1 avector00_reg_5__5_ ( .D(n21543), .CK(clk), .QN(n18547) );
  DFF_X1 avector00_reg_5__6_ ( .D(n21542), .CK(clk), .QN(n18510) );
  DFF_X1 avector00_reg_5__7_ ( .D(n21541), .CK(clk), .QN(n18473) );
  DFF_X1 avector00_reg_5__8_ ( .D(n21540), .CK(clk), .QN(n18436) );
  DFF_X1 avector00_reg_5__9_ ( .D(n21539), .CK(clk), .QN(n18399) );
  DFF_X1 avector00_reg_5__10_ ( .D(n21538), .CK(clk), .QN(n18362) );
  DFF_X1 avector00_reg_5__11_ ( .D(n21537), .CK(clk), .QN(n18325) );
  DFF_X1 avector00_reg_5__12_ ( .D(n21536), .CK(clk), .QN(n18288) );
  DFF_X1 avector00_reg_5__13_ ( .D(n21535), .CK(clk), .QN(n18251) );
  DFF_X1 avector00_reg_5__14_ ( .D(n21534), .CK(clk), .QN(n18214) );
  DFF_X1 avector00_reg_5__15_ ( .D(n21533), .CK(clk), .QN(n18177) );
  DFF_X1 avector30_reg_5__0_ ( .D(n21484), .CK(clk), .QN(n16956) );
  DFF_X1 avector30_reg_5__1_ ( .D(n21483), .CK(clk), .QN(n16919) );
  DFF_X1 avector30_reg_5__2_ ( .D(n21482), .CK(clk), .QN(n16882) );
  DFF_X1 avector30_reg_5__3_ ( .D(n21481), .CK(clk), .QN(n16845) );
  DFF_X1 avector30_reg_5__4_ ( .D(n21480), .CK(clk), .QN(n16808) );
  DFF_X1 avector30_reg_5__5_ ( .D(n21479), .CK(clk), .QN(n16771) );
  DFF_X1 avector30_reg_5__6_ ( .D(n21478), .CK(clk), .QN(n16734) );
  DFF_X1 avector30_reg_5__7_ ( .D(n21477), .CK(clk), .QN(n16697) );
  DFF_X1 avector30_reg_5__8_ ( .D(n21476), .CK(clk), .QN(n16660) );
  DFF_X1 avector30_reg_5__9_ ( .D(n21475), .CK(clk), .QN(n16623) );
  DFF_X1 avector30_reg_5__10_ ( .D(n21474), .CK(clk), .QN(n16586) );
  DFF_X1 avector30_reg_5__11_ ( .D(n21473), .CK(clk), .QN(n16549) );
  DFF_X1 avector30_reg_5__12_ ( .D(n21472), .CK(clk), .QN(n16512) );
  DFF_X1 avector30_reg_5__13_ ( .D(n21471), .CK(clk), .QN(n16475) );
  DFF_X1 avector30_reg_5__14_ ( .D(n21470), .CK(clk), .QN(n16438) );
  DFF_X1 avector30_reg_5__15_ ( .D(n21469), .CK(clk), .QN(n16401) );
  DFF_X1 avector23_reg_3__0_ ( .D(n22348), .CK(clk), .QN(n17552) );
  DFF_X1 avector23_reg_3__1_ ( .D(n22347), .CK(clk), .QN(n17515) );
  DFF_X1 avector23_reg_3__2_ ( .D(n22346), .CK(clk), .QN(n17478) );
  DFF_X1 avector23_reg_3__3_ ( .D(n22345), .CK(clk), .QN(n17441) );
  DFF_X1 avector23_reg_3__4_ ( .D(n22344), .CK(clk), .QN(n17404) );
  DFF_X1 avector23_reg_3__5_ ( .D(n22343), .CK(clk), .QN(n17367) );
  DFF_X1 avector23_reg_3__6_ ( .D(n22342), .CK(clk), .QN(n17330) );
  DFF_X1 avector23_reg_3__7_ ( .D(n22341), .CK(clk), .QN(n17293) );
  DFF_X1 avector23_reg_3__8_ ( .D(n22340), .CK(clk), .QN(n17256) );
  DFF_X1 avector23_reg_3__9_ ( .D(n22339), .CK(clk), .QN(n17219) );
  DFF_X1 avector23_reg_3__10_ ( .D(n22338), .CK(clk), .QN(n17182) );
  DFF_X1 avector23_reg_3__11_ ( .D(n22337), .CK(clk), .QN(n17145) );
  DFF_X1 avector23_reg_3__12_ ( .D(n22336), .CK(clk), .QN(n17108) );
  DFF_X1 avector23_reg_3__13_ ( .D(n22335), .CK(clk), .QN(n17071) );
  DFF_X1 avector23_reg_3__14_ ( .D(n22334), .CK(clk), .QN(n17034) );
  DFF_X1 avector23_reg_3__15_ ( .D(n22333), .CK(clk), .QN(n16997) );
  DFF_X1 avector13_reg_3__0_ ( .D(n22284), .CK(clk), .QN(n18144) );
  DFF_X1 avector13_reg_3__1_ ( .D(n22283), .CK(clk), .QN(n18107) );
  DFF_X1 avector13_reg_3__2_ ( .D(n22282), .CK(clk), .QN(n18070) );
  DFF_X1 avector13_reg_3__3_ ( .D(n22281), .CK(clk), .QN(n18033) );
  DFF_X1 avector13_reg_3__4_ ( .D(n22280), .CK(clk), .QN(n17996) );
  DFF_X1 avector13_reg_3__5_ ( .D(n22279), .CK(clk), .QN(n17959) );
  DFF_X1 avector13_reg_3__6_ ( .D(n22278), .CK(clk), .QN(n17922) );
  DFF_X1 avector13_reg_3__7_ ( .D(n22277), .CK(clk), .QN(n17885) );
  DFF_X1 avector13_reg_3__8_ ( .D(n22276), .CK(clk), .QN(n17848) );
  DFF_X1 avector13_reg_3__9_ ( .D(n22275), .CK(clk), .QN(n17811) );
  DFF_X1 avector13_reg_3__10_ ( .D(n22274), .CK(clk), .QN(n17774) );
  DFF_X1 avector13_reg_3__11_ ( .D(n22273), .CK(clk), .QN(n17737) );
  DFF_X1 avector13_reg_3__12_ ( .D(n22272), .CK(clk), .QN(n17700) );
  DFF_X1 avector13_reg_3__13_ ( .D(n22271), .CK(clk), .QN(n17663) );
  DFF_X1 avector13_reg_3__14_ ( .D(n22270), .CK(clk), .QN(n17626) );
  DFF_X1 avector13_reg_3__15_ ( .D(n22269), .CK(clk), .QN(n17589) );
  DFF_X1 avector03_reg_3__0_ ( .D(n22220), .CK(clk), .QN(n18736) );
  DFF_X1 avector03_reg_3__1_ ( .D(n22219), .CK(clk), .QN(n18699) );
  DFF_X1 avector03_reg_3__2_ ( .D(n22218), .CK(clk), .QN(n18662) );
  DFF_X1 avector03_reg_3__3_ ( .D(n22217), .CK(clk), .QN(n18625) );
  DFF_X1 avector03_reg_3__4_ ( .D(n22216), .CK(clk), .QN(n18588) );
  DFF_X1 avector03_reg_3__5_ ( .D(n22215), .CK(clk), .QN(n18551) );
  DFF_X1 avector03_reg_3__6_ ( .D(n22214), .CK(clk), .QN(n18514) );
  DFF_X1 avector03_reg_3__7_ ( .D(n22213), .CK(clk), .QN(n18477) );
  DFF_X1 avector03_reg_3__8_ ( .D(n22212), .CK(clk), .QN(n18440) );
  DFF_X1 avector03_reg_3__9_ ( .D(n22211), .CK(clk), .QN(n18403) );
  DFF_X1 avector03_reg_3__10_ ( .D(n22210), .CK(clk), .QN(n18366) );
  DFF_X1 avector03_reg_3__11_ ( .D(n22209), .CK(clk), .QN(n18329) );
  DFF_X1 avector03_reg_3__12_ ( .D(n22208), .CK(clk), .QN(n18292) );
  DFF_X1 avector03_reg_3__13_ ( .D(n22207), .CK(clk), .QN(n18255) );
  DFF_X1 avector03_reg_3__14_ ( .D(n22206), .CK(clk), .QN(n18218) );
  DFF_X1 avector03_reg_3__15_ ( .D(n22205), .CK(clk), .QN(n18181) );
  DFF_X1 avector33_reg_3__0_ ( .D(n21116), .CK(clk), .QN(n16960) );
  DFF_X1 avector33_reg_3__1_ ( .D(n21115), .CK(clk), .QN(n16923) );
  DFF_X1 avector33_reg_3__2_ ( .D(n21114), .CK(clk), .QN(n16886) );
  DFF_X1 avector33_reg_3__3_ ( .D(n21113), .CK(clk), .QN(n16849) );
  DFF_X1 avector33_reg_3__4_ ( .D(n21112), .CK(clk), .QN(n16812) );
  DFF_X1 avector33_reg_3__5_ ( .D(n21111), .CK(clk), .QN(n16775) );
  DFF_X1 avector33_reg_3__6_ ( .D(n21110), .CK(clk), .QN(n16738) );
  DFF_X1 avector33_reg_3__7_ ( .D(n21109), .CK(clk), .QN(n16701) );
  DFF_X1 avector33_reg_3__8_ ( .D(n21108), .CK(clk), .QN(n16664) );
  DFF_X1 avector33_reg_3__9_ ( .D(n21107), .CK(clk), .QN(n16627) );
  DFF_X1 avector33_reg_3__10_ ( .D(n21106), .CK(clk), .QN(n16590) );
  DFF_X1 avector33_reg_3__11_ ( .D(n21105), .CK(clk), .QN(n16553) );
  DFF_X1 avector33_reg_3__12_ ( .D(n21104), .CK(clk), .QN(n16516) );
  DFF_X1 avector33_reg_3__13_ ( .D(n21103), .CK(clk), .QN(n16479) );
  DFF_X1 avector33_reg_3__14_ ( .D(n21102), .CK(clk), .QN(n16442) );
  DFF_X1 avector33_reg_3__15_ ( .D(n21101), .CK(clk), .QN(n16405) );
  DFF_X1 avector22_reg_3__0_ ( .D(n22156), .CK(clk), .QN(n17525) );
  DFF_X1 avector22_reg_3__1_ ( .D(n22155), .CK(clk), .QN(n17488) );
  DFF_X1 avector22_reg_3__2_ ( .D(n22154), .CK(clk), .QN(n17451) );
  DFF_X1 avector22_reg_3__3_ ( .D(n22153), .CK(clk), .QN(n17414) );
  DFF_X1 avector22_reg_3__4_ ( .D(n22152), .CK(clk), .QN(n17377) );
  DFF_X1 avector22_reg_3__5_ ( .D(n22151), .CK(clk), .QN(n17340) );
  DFF_X1 avector22_reg_3__6_ ( .D(n22150), .CK(clk), .QN(n17303) );
  DFF_X1 avector22_reg_3__7_ ( .D(n22149), .CK(clk), .QN(n17266) );
  DFF_X1 avector22_reg_3__8_ ( .D(n22148), .CK(clk), .QN(n17229) );
  DFF_X1 avector22_reg_3__9_ ( .D(n22147), .CK(clk), .QN(n17192) );
  DFF_X1 avector22_reg_3__10_ ( .D(n22146), .CK(clk), .QN(n17155) );
  DFF_X1 avector22_reg_3__11_ ( .D(n22145), .CK(clk), .QN(n17118) );
  DFF_X1 avector22_reg_3__12_ ( .D(n22144), .CK(clk), .QN(n17081) );
  DFF_X1 avector22_reg_3__13_ ( .D(n22143), .CK(clk), .QN(n17044) );
  DFF_X1 avector22_reg_3__14_ ( .D(n22142), .CK(clk), .QN(n17007) );
  DFF_X1 avector22_reg_3__15_ ( .D(n22141), .CK(clk), .QN(n16970) );
  DFF_X1 avector12_reg_3__0_ ( .D(n22092), .CK(clk), .QN(n18117) );
  DFF_X1 avector12_reg_3__1_ ( .D(n22091), .CK(clk), .QN(n18080) );
  DFF_X1 avector12_reg_3__2_ ( .D(n22090), .CK(clk), .QN(n18043) );
  DFF_X1 avector12_reg_3__3_ ( .D(n22089), .CK(clk), .QN(n18006) );
  DFF_X1 avector12_reg_3__4_ ( .D(n22088), .CK(clk), .QN(n17969) );
  DFF_X1 avector12_reg_3__5_ ( .D(n22087), .CK(clk), .QN(n17932) );
  DFF_X1 avector12_reg_3__6_ ( .D(n22086), .CK(clk), .QN(n17895) );
  DFF_X1 avector12_reg_3__7_ ( .D(n22085), .CK(clk), .QN(n17858) );
  DFF_X1 avector12_reg_3__8_ ( .D(n22084), .CK(clk), .QN(n17821) );
  DFF_X1 avector12_reg_3__9_ ( .D(n22083), .CK(clk), .QN(n17784) );
  DFF_X1 avector12_reg_3__10_ ( .D(n22082), .CK(clk), .QN(n17747) );
  DFF_X1 avector12_reg_3__11_ ( .D(n22081), .CK(clk), .QN(n17710) );
  DFF_X1 avector12_reg_3__12_ ( .D(n22080), .CK(clk), .QN(n17673) );
  DFF_X1 avector12_reg_3__13_ ( .D(n22079), .CK(clk), .QN(n17636) );
  DFF_X1 avector12_reg_3__14_ ( .D(n22078), .CK(clk), .QN(n17599) );
  DFF_X1 avector12_reg_3__15_ ( .D(n22077), .CK(clk), .QN(n17562) );
  DFF_X1 avector02_reg_3__0_ ( .D(n22028), .CK(clk), .QN(n18709) );
  DFF_X1 avector02_reg_3__1_ ( .D(n22027), .CK(clk), .QN(n18672) );
  DFF_X1 avector02_reg_3__2_ ( .D(n22026), .CK(clk), .QN(n18635) );
  DFF_X1 avector02_reg_3__3_ ( .D(n22025), .CK(clk), .QN(n18598) );
  DFF_X1 avector02_reg_3__4_ ( .D(n22024), .CK(clk), .QN(n18561) );
  DFF_X1 avector02_reg_3__5_ ( .D(n22023), .CK(clk), .QN(n18524) );
  DFF_X1 avector02_reg_3__6_ ( .D(n22022), .CK(clk), .QN(n18487) );
  DFF_X1 avector02_reg_3__7_ ( .D(n22021), .CK(clk), .QN(n18450) );
  DFF_X1 avector02_reg_3__8_ ( .D(n22020), .CK(clk), .QN(n18413) );
  DFF_X1 avector02_reg_3__9_ ( .D(n22019), .CK(clk), .QN(n18376) );
  DFF_X1 avector02_reg_3__10_ ( .D(n22018), .CK(clk), .QN(n18339) );
  DFF_X1 avector02_reg_3__11_ ( .D(n22017), .CK(clk), .QN(n18302) );
  DFF_X1 avector02_reg_3__12_ ( .D(n22016), .CK(clk), .QN(n18265) );
  DFF_X1 avector02_reg_3__13_ ( .D(n22015), .CK(clk), .QN(n18228) );
  DFF_X1 avector02_reg_3__14_ ( .D(n22014), .CK(clk), .QN(n18191) );
  DFF_X1 avector02_reg_3__15_ ( .D(n22013), .CK(clk), .QN(n18154) );
  DFF_X1 avector32_reg_3__0_ ( .D(n21964), .CK(clk), .QN(n16933) );
  DFF_X1 avector32_reg_3__1_ ( .D(n21963), .CK(clk), .QN(n16896) );
  DFF_X1 avector32_reg_3__2_ ( .D(n21962), .CK(clk), .QN(n16859) );
  DFF_X1 avector32_reg_3__3_ ( .D(n21961), .CK(clk), .QN(n16822) );
  DFF_X1 avector32_reg_3__4_ ( .D(n21960), .CK(clk), .QN(n16785) );
  DFF_X1 avector32_reg_3__5_ ( .D(n21959), .CK(clk), .QN(n16748) );
  DFF_X1 avector32_reg_3__6_ ( .D(n21958), .CK(clk), .QN(n16711) );
  DFF_X1 avector32_reg_3__7_ ( .D(n21957), .CK(clk), .QN(n16674) );
  DFF_X1 avector32_reg_3__8_ ( .D(n21956), .CK(clk), .QN(n16637) );
  DFF_X1 avector32_reg_3__9_ ( .D(n21955), .CK(clk), .QN(n16600) );
  DFF_X1 avector32_reg_3__10_ ( .D(n21954), .CK(clk), .QN(n16563) );
  DFF_X1 avector32_reg_3__11_ ( .D(n21953), .CK(clk), .QN(n16526) );
  DFF_X1 avector32_reg_3__12_ ( .D(n21952), .CK(clk), .QN(n16489) );
  DFF_X1 avector32_reg_3__13_ ( .D(n21951), .CK(clk), .QN(n16452) );
  DFF_X1 avector32_reg_3__14_ ( .D(n21950), .CK(clk), .QN(n16415) );
  DFF_X1 avector32_reg_3__15_ ( .D(n21949), .CK(clk), .QN(n16378) );
  DFF_X1 avector21_reg_3__0_ ( .D(n21900), .CK(clk), .Q(n25470), .QN(n17534)
         );
  DFF_X1 avector21_reg_3__1_ ( .D(n21899), .CK(clk), .Q(n25467), .QN(n17497)
         );
  DFF_X1 avector21_reg_3__2_ ( .D(n21898), .CK(clk), .Q(n25464), .QN(n17460)
         );
  DFF_X1 avector21_reg_3__3_ ( .D(n21897), .CK(clk), .Q(n25461), .QN(n17423)
         );
  DFF_X1 avector21_reg_3__4_ ( .D(n21896), .CK(clk), .Q(n25458), .QN(n17386)
         );
  DFF_X1 avector21_reg_3__5_ ( .D(n21895), .CK(clk), .Q(n25455), .QN(n17349)
         );
  DFF_X1 avector21_reg_3__6_ ( .D(n21894), .CK(clk), .Q(n25452), .QN(n17312)
         );
  DFF_X1 avector21_reg_3__7_ ( .D(n21893), .CK(clk), .Q(n25449), .QN(n17275)
         );
  DFF_X1 avector21_reg_3__8_ ( .D(n21892), .CK(clk), .Q(n25446), .QN(n17238)
         );
  DFF_X1 avector21_reg_3__9_ ( .D(n21891), .CK(clk), .Q(n25443), .QN(n17201)
         );
  DFF_X1 avector21_reg_3__10_ ( .D(n21890), .CK(clk), .Q(n25440), .QN(n17164)
         );
  DFF_X1 avector21_reg_3__11_ ( .D(n21889), .CK(clk), .Q(n25437), .QN(n17127)
         );
  DFF_X1 avector21_reg_3__12_ ( .D(n21888), .CK(clk), .Q(n25149), .QN(n17090)
         );
  DFF_X1 avector21_reg_3__13_ ( .D(n21887), .CK(clk), .Q(n25146), .QN(n17053)
         );
  DFF_X1 avector21_reg_3__14_ ( .D(n21886), .CK(clk), .Q(n25143), .QN(n17016)
         );
  DFF_X1 avector21_reg_3__15_ ( .D(n21885), .CK(clk), .Q(n25140), .QN(n16979)
         );
  DFF_X1 avector11_reg_3__0_ ( .D(n21836), .CK(clk), .Q(n25510), .QN(n18126)
         );
  DFF_X1 avector11_reg_3__1_ ( .D(n21835), .CK(clk), .Q(n25507), .QN(n18089)
         );
  DFF_X1 avector11_reg_3__2_ ( .D(n21834), .CK(clk), .Q(n25504), .QN(n18052)
         );
  DFF_X1 avector11_reg_3__3_ ( .D(n21833), .CK(clk), .Q(n25501), .QN(n18015)
         );
  DFF_X1 avector11_reg_3__4_ ( .D(n21832), .CK(clk), .Q(n25498), .QN(n17978)
         );
  DFF_X1 avector11_reg_3__5_ ( .D(n21831), .CK(clk), .Q(n25495), .QN(n17941)
         );
  DFF_X1 avector11_reg_3__6_ ( .D(n21830), .CK(clk), .Q(n25492), .QN(n17904)
         );
  DFF_X1 avector11_reg_3__7_ ( .D(n21829), .CK(clk), .Q(n25489), .QN(n17867)
         );
  DFF_X1 avector11_reg_3__8_ ( .D(n21828), .CK(clk), .Q(n25486), .QN(n17830)
         );
  DFF_X1 avector11_reg_3__9_ ( .D(n21827), .CK(clk), .Q(n25483), .QN(n17793)
         );
  DFF_X1 avector11_reg_3__10_ ( .D(n21826), .CK(clk), .Q(n25480), .QN(n17756)
         );
  DFF_X1 avector11_reg_3__11_ ( .D(n21825), .CK(clk), .Q(n25477), .QN(n17719)
         );
  DFF_X1 avector11_reg_3__12_ ( .D(n21824), .CK(clk), .Q(n25173), .QN(n17682)
         );
  DFF_X1 avector11_reg_3__13_ ( .D(n21823), .CK(clk), .Q(n25170), .QN(n17645)
         );
  DFF_X1 avector11_reg_3__14_ ( .D(n21822), .CK(clk), .Q(n25167), .QN(n17608)
         );
  DFF_X1 avector11_reg_3__15_ ( .D(n21821), .CK(clk), .Q(n25164), .QN(n17571)
         );
  DFF_X1 avector01_reg_3__0_ ( .D(n21772), .CK(clk), .Q(n25550), .QN(n18718)
         );
  DFF_X1 avector01_reg_3__1_ ( .D(n21771), .CK(clk), .Q(n25547), .QN(n18681)
         );
  DFF_X1 avector01_reg_3__2_ ( .D(n21770), .CK(clk), .Q(n25544), .QN(n18644)
         );
  DFF_X1 avector01_reg_3__3_ ( .D(n21769), .CK(clk), .Q(n25541), .QN(n18607)
         );
  DFF_X1 avector01_reg_3__4_ ( .D(n21768), .CK(clk), .Q(n25538), .QN(n18570)
         );
  DFF_X1 avector01_reg_3__5_ ( .D(n21767), .CK(clk), .Q(n25535), .QN(n18533)
         );
  DFF_X1 avector01_reg_3__6_ ( .D(n21766), .CK(clk), .Q(n25532), .QN(n18496)
         );
  DFF_X1 avector01_reg_3__7_ ( .D(n21765), .CK(clk), .Q(n25529), .QN(n18459)
         );
  DFF_X1 avector01_reg_3__8_ ( .D(n21764), .CK(clk), .Q(n25526), .QN(n18422)
         );
  DFF_X1 avector01_reg_3__9_ ( .D(n21763), .CK(clk), .Q(n25523), .QN(n18385)
         );
  DFF_X1 avector01_reg_3__10_ ( .D(n21762), .CK(clk), .Q(n25520), .QN(n18348)
         );
  DFF_X1 avector01_reg_3__11_ ( .D(n21761), .CK(clk), .Q(n25517), .QN(n18311)
         );
  DFF_X1 avector01_reg_3__12_ ( .D(n21760), .CK(clk), .Q(n25197), .QN(n18274)
         );
  DFF_X1 avector01_reg_3__13_ ( .D(n21759), .CK(clk), .Q(n25194), .QN(n18237)
         );
  DFF_X1 avector01_reg_3__14_ ( .D(n21758), .CK(clk), .Q(n25191), .QN(n18200)
         );
  DFF_X1 avector01_reg_3__15_ ( .D(n21757), .CK(clk), .Q(n25188), .QN(n18163)
         );
  DFF_X1 avector31_reg_3__0_ ( .D(n21708), .CK(clk), .Q(n25430), .QN(n16942)
         );
  DFF_X1 avector31_reg_3__1_ ( .D(n21707), .CK(clk), .Q(n25427), .QN(n16905)
         );
  DFF_X1 avector31_reg_3__2_ ( .D(n21706), .CK(clk), .Q(n25423), .QN(n16868)
         );
  DFF_X1 avector31_reg_3__3_ ( .D(n21705), .CK(clk), .Q(n25420), .QN(n16831)
         );
  DFF_X1 avector31_reg_3__4_ ( .D(n21704), .CK(clk), .Q(n25417), .QN(n16794)
         );
  DFF_X1 avector31_reg_3__5_ ( .D(n21703), .CK(clk), .Q(n25414), .QN(n16757)
         );
  DFF_X1 avector31_reg_3__6_ ( .D(n21702), .CK(clk), .Q(n25133), .QN(n16720)
         );
  DFF_X1 avector31_reg_3__7_ ( .D(n21701), .CK(clk), .Q(n25130), .QN(n16683)
         );
  DFF_X1 avector31_reg_3__8_ ( .D(n21700), .CK(clk), .Q(n25127), .QN(n16646)
         );
  DFF_X1 avector31_reg_3__9_ ( .D(n21699), .CK(clk), .Q(n25124), .QN(n16609)
         );
  DFF_X1 avector31_reg_3__10_ ( .D(n21698), .CK(clk), .Q(n25121), .QN(n16572)
         );
  DFF_X1 avector31_reg_3__11_ ( .D(n21697), .CK(clk), .Q(n25118), .QN(n16535)
         );
  DFF_X1 avector31_reg_3__12_ ( .D(n21696), .CK(clk), .Q(n25115), .QN(n16498)
         );
  DFF_X1 avector31_reg_3__13_ ( .D(n21695), .CK(clk), .Q(n25112), .QN(n16461)
         );
  DFF_X1 avector31_reg_3__14_ ( .D(n21694), .CK(clk), .Q(n25109), .QN(n16424)
         );
  DFF_X1 avector31_reg_3__15_ ( .D(n21693), .CK(clk), .Q(n25106), .QN(n16387)
         );
  DFF_X1 avector20_reg_3__0_ ( .D(n21644), .CK(clk), .Q(n25003), .QN(n17543)
         );
  DFF_X1 avector20_reg_3__1_ ( .D(n21643), .CK(clk), .Q(n25001), .QN(n17506)
         );
  DFF_X1 avector20_reg_3__2_ ( .D(n21642), .CK(clk), .Q(n24999), .QN(n17469)
         );
  DFF_X1 avector20_reg_3__3_ ( .D(n21641), .CK(clk), .Q(n24997), .QN(n17432)
         );
  DFF_X1 avector20_reg_3__4_ ( .D(n21640), .CK(clk), .Q(n24995), .QN(n17395)
         );
  DFF_X1 avector20_reg_3__5_ ( .D(n21639), .CK(clk), .Q(n24993), .QN(n17358)
         );
  DFF_X1 avector20_reg_3__6_ ( .D(n21638), .CK(clk), .Q(n24991), .QN(n17321)
         );
  DFF_X1 avector20_reg_3__7_ ( .D(n21637), .CK(clk), .Q(n24989), .QN(n17284)
         );
  DFF_X1 avector20_reg_3__8_ ( .D(n21636), .CK(clk), .Q(n24987), .QN(n17247)
         );
  DFF_X1 avector20_reg_3__9_ ( .D(n21635), .CK(clk), .Q(n24985), .QN(n17210)
         );
  DFF_X1 avector20_reg_3__10_ ( .D(n21634), .CK(clk), .Q(n24983), .QN(n17173)
         );
  DFF_X1 avector20_reg_3__11_ ( .D(n21633), .CK(clk), .Q(n24981), .QN(n17136)
         );
  DFF_X1 avector20_reg_3__12_ ( .D(n21632), .CK(clk), .Q(n25636), .QN(n17099)
         );
  DFF_X1 avector20_reg_3__13_ ( .D(n21631), .CK(clk), .Q(n25633), .QN(n17062)
         );
  DFF_X1 avector20_reg_3__14_ ( .D(n21630), .CK(clk), .Q(n25630), .QN(n17025)
         );
  DFF_X1 avector20_reg_3__15_ ( .D(n21629), .CK(clk), .Q(n25627), .QN(n16988)
         );
  DFF_X1 avector10_reg_3__0_ ( .D(n21580), .CK(clk), .Q(n25027), .QN(n18135)
         );
  DFF_X1 avector10_reg_3__1_ ( .D(n21579), .CK(clk), .Q(n25025), .QN(n18098)
         );
  DFF_X1 avector10_reg_3__2_ ( .D(n21578), .CK(clk), .Q(n25023), .QN(n18061)
         );
  DFF_X1 avector10_reg_3__3_ ( .D(n21577), .CK(clk), .Q(n25021), .QN(n18024)
         );
  DFF_X1 avector10_reg_3__4_ ( .D(n21576), .CK(clk), .Q(n25019), .QN(n17987)
         );
  DFF_X1 avector10_reg_3__5_ ( .D(n21575), .CK(clk), .Q(n25017), .QN(n17950)
         );
  DFF_X1 avector10_reg_3__6_ ( .D(n21574), .CK(clk), .Q(n25015), .QN(n17913)
         );
  DFF_X1 avector10_reg_3__7_ ( .D(n21573), .CK(clk), .Q(n25013), .QN(n17876)
         );
  DFF_X1 avector10_reg_3__8_ ( .D(n21572), .CK(clk), .Q(n25011), .QN(n17839)
         );
  DFF_X1 avector10_reg_3__9_ ( .D(n21571), .CK(clk), .Q(n25009), .QN(n17802)
         );
  DFF_X1 avector10_reg_3__10_ ( .D(n21570), .CK(clk), .Q(n25007), .QN(n17765)
         );
  DFF_X1 avector10_reg_3__11_ ( .D(n21569), .CK(clk), .Q(n25005), .QN(n17728)
         );
  DFF_X1 avector10_reg_3__12_ ( .D(n21568), .CK(clk), .Q(n25660), .QN(n17691)
         );
  DFF_X1 avector10_reg_3__13_ ( .D(n21567), .CK(clk), .Q(n25657), .QN(n17654)
         );
  DFF_X1 avector10_reg_3__14_ ( .D(n21566), .CK(clk), .Q(n25654), .QN(n17617)
         );
  DFF_X1 avector10_reg_3__15_ ( .D(n21565), .CK(clk), .Q(n25651), .QN(n17580)
         );
  DFF_X1 avector00_reg_3__0_ ( .D(n21516), .CK(clk), .Q(n25051), .QN(n18727)
         );
  DFF_X1 avector00_reg_3__1_ ( .D(n21515), .CK(clk), .Q(n25049), .QN(n18690)
         );
  DFF_X1 avector00_reg_3__2_ ( .D(n21514), .CK(clk), .Q(n25047), .QN(n18653)
         );
  DFF_X1 avector00_reg_3__3_ ( .D(n21513), .CK(clk), .Q(n25045), .QN(n18616)
         );
  DFF_X1 avector00_reg_3__4_ ( .D(n21512), .CK(clk), .Q(n25043), .QN(n18579)
         );
  DFF_X1 avector00_reg_3__5_ ( .D(n21511), .CK(clk), .Q(n25041), .QN(n18542)
         );
  DFF_X1 avector00_reg_3__6_ ( .D(n21510), .CK(clk), .Q(n25039), .QN(n18505)
         );
  DFF_X1 avector00_reg_3__7_ ( .D(n21509), .CK(clk), .Q(n25037), .QN(n18468)
         );
  DFF_X1 avector00_reg_3__8_ ( .D(n21508), .CK(clk), .Q(n25035), .QN(n18431)
         );
  DFF_X1 avector00_reg_3__9_ ( .D(n21507), .CK(clk), .Q(n25033), .QN(n18394)
         );
  DFF_X1 avector00_reg_3__10_ ( .D(n21506), .CK(clk), .Q(n25031), .QN(n18357)
         );
  DFF_X1 avector00_reg_3__11_ ( .D(n21505), .CK(clk), .Q(n25029), .QN(n18320)
         );
  DFF_X1 avector00_reg_3__12_ ( .D(n21504), .CK(clk), .Q(n25684), .QN(n18283)
         );
  DFF_X1 avector00_reg_3__13_ ( .D(n21503), .CK(clk), .Q(n25681), .QN(n18246)
         );
  DFF_X1 avector00_reg_3__14_ ( .D(n21502), .CK(clk), .Q(n25678), .QN(n18209)
         );
  DFF_X1 avector00_reg_3__15_ ( .D(n21501), .CK(clk), .Q(n25675), .QN(n18172)
         );
  DFF_X1 avector30_reg_3__0_ ( .D(n21452), .CK(clk), .Q(n24979), .QN(n16951)
         );
  DFF_X1 avector30_reg_3__1_ ( .D(n21451), .CK(clk), .Q(n24977), .QN(n16914)
         );
  DFF_X1 avector30_reg_3__2_ ( .D(n21450), .CK(clk), .Q(n24974), .QN(n16877)
         );
  DFF_X1 avector30_reg_3__3_ ( .D(n21449), .CK(clk), .Q(n24972), .QN(n16840)
         );
  DFF_X1 avector30_reg_3__4_ ( .D(n21448), .CK(clk), .Q(n24970), .QN(n16803)
         );
  DFF_X1 avector30_reg_3__5_ ( .D(n21447), .CK(clk), .Q(n24968), .QN(n16766)
         );
  DFF_X1 avector30_reg_3__6_ ( .D(n21446), .CK(clk), .Q(n25620), .QN(n16729)
         );
  DFF_X1 avector30_reg_3__7_ ( .D(n21445), .CK(clk), .Q(n25617), .QN(n16692)
         );
  DFF_X1 avector30_reg_3__8_ ( .D(n21444), .CK(clk), .Q(n25614), .QN(n16655)
         );
  DFF_X1 avector30_reg_3__9_ ( .D(n21443), .CK(clk), .Q(n25611), .QN(n16618)
         );
  DFF_X1 avector30_reg_3__10_ ( .D(n21442), .CK(clk), .Q(n25608), .QN(n16581)
         );
  DFF_X1 avector30_reg_3__11_ ( .D(n21441), .CK(clk), .Q(n25605), .QN(n16544)
         );
  DFF_X1 avector30_reg_3__12_ ( .D(n21440), .CK(clk), .Q(n25602), .QN(n16507)
         );
  DFF_X1 avector30_reg_3__13_ ( .D(n21439), .CK(clk), .Q(n25599), .QN(n16470)
         );
  DFF_X1 avector30_reg_3__14_ ( .D(n21438), .CK(clk), .Q(n25596), .QN(n16433)
         );
  DFF_X1 avector30_reg_3__15_ ( .D(n21437), .CK(clk), .Q(n25593), .QN(n16396)
         );
  DFF_X1 avector23_reg_2__0_ ( .D(n22332), .CK(clk), .QN(n17551) );
  DFF_X1 avector23_reg_2__1_ ( .D(n22331), .CK(clk), .QN(n17514) );
  DFF_X1 avector23_reg_2__2_ ( .D(n22330), .CK(clk), .QN(n17477) );
  DFF_X1 avector23_reg_2__3_ ( .D(n22329), .CK(clk), .QN(n17440) );
  DFF_X1 avector23_reg_2__4_ ( .D(n22328), .CK(clk), .QN(n17403) );
  DFF_X1 avector23_reg_2__5_ ( .D(n22327), .CK(clk), .QN(n17366) );
  DFF_X1 avector23_reg_2__6_ ( .D(n22326), .CK(clk), .QN(n17329) );
  DFF_X1 avector23_reg_2__7_ ( .D(n22325), .CK(clk), .QN(n17292) );
  DFF_X1 avector23_reg_2__8_ ( .D(n22324), .CK(clk), .QN(n17255) );
  DFF_X1 avector23_reg_2__9_ ( .D(n22323), .CK(clk), .QN(n17218) );
  DFF_X1 avector23_reg_2__10_ ( .D(n22322), .CK(clk), .QN(n17181) );
  DFF_X1 avector23_reg_2__11_ ( .D(n22321), .CK(clk), .QN(n17144) );
  DFF_X1 avector23_reg_2__12_ ( .D(n22320), .CK(clk), .QN(n17107) );
  DFF_X1 avector23_reg_2__13_ ( .D(n22319), .CK(clk), .QN(n17070) );
  DFF_X1 avector23_reg_2__14_ ( .D(n22318), .CK(clk), .QN(n17033) );
  DFF_X1 avector23_reg_2__15_ ( .D(n22317), .CK(clk), .QN(n16996) );
  DFF_X1 avector13_reg_2__0_ ( .D(n22268), .CK(clk), .QN(n18143) );
  DFF_X1 avector13_reg_2__1_ ( .D(n22267), .CK(clk), .QN(n18106) );
  DFF_X1 avector13_reg_2__2_ ( .D(n22266), .CK(clk), .QN(n18069) );
  DFF_X1 avector13_reg_2__3_ ( .D(n22265), .CK(clk), .QN(n18032) );
  DFF_X1 avector13_reg_2__4_ ( .D(n22264), .CK(clk), .QN(n17995) );
  DFF_X1 avector13_reg_2__5_ ( .D(n22263), .CK(clk), .QN(n17958) );
  DFF_X1 avector13_reg_2__6_ ( .D(n22262), .CK(clk), .QN(n17921) );
  DFF_X1 avector13_reg_2__7_ ( .D(n22261), .CK(clk), .QN(n17884) );
  DFF_X1 avector13_reg_2__8_ ( .D(n22260), .CK(clk), .QN(n17847) );
  DFF_X1 avector13_reg_2__9_ ( .D(n22259), .CK(clk), .QN(n17810) );
  DFF_X1 avector13_reg_2__10_ ( .D(n22258), .CK(clk), .QN(n17773) );
  DFF_X1 avector13_reg_2__11_ ( .D(n22257), .CK(clk), .QN(n17736) );
  DFF_X1 avector13_reg_2__12_ ( .D(n22256), .CK(clk), .QN(n17699) );
  DFF_X1 avector13_reg_2__13_ ( .D(n22255), .CK(clk), .QN(n17662) );
  DFF_X1 avector13_reg_2__14_ ( .D(n22254), .CK(clk), .QN(n17625) );
  DFF_X1 avector13_reg_2__15_ ( .D(n22253), .CK(clk), .QN(n17588) );
  DFF_X1 avector03_reg_2__0_ ( .D(n22204), .CK(clk), .QN(n18735) );
  DFF_X1 avector03_reg_2__1_ ( .D(n22203), .CK(clk), .QN(n18698) );
  DFF_X1 avector03_reg_2__2_ ( .D(n22202), .CK(clk), .QN(n18661) );
  DFF_X1 avector03_reg_2__3_ ( .D(n22201), .CK(clk), .QN(n18624) );
  DFF_X1 avector03_reg_2__4_ ( .D(n22200), .CK(clk), .QN(n18587) );
  DFF_X1 avector03_reg_2__5_ ( .D(n22199), .CK(clk), .QN(n18550) );
  DFF_X1 avector03_reg_2__6_ ( .D(n22198), .CK(clk), .QN(n18513) );
  DFF_X1 avector03_reg_2__7_ ( .D(n22197), .CK(clk), .QN(n18476) );
  DFF_X1 avector03_reg_2__8_ ( .D(n22196), .CK(clk), .QN(n18439) );
  DFF_X1 avector03_reg_2__9_ ( .D(n22195), .CK(clk), .QN(n18402) );
  DFF_X1 avector03_reg_2__10_ ( .D(n22194), .CK(clk), .QN(n18365) );
  DFF_X1 avector03_reg_2__11_ ( .D(n22193), .CK(clk), .QN(n18328) );
  DFF_X1 avector03_reg_2__12_ ( .D(n22192), .CK(clk), .QN(n18291) );
  DFF_X1 avector03_reg_2__13_ ( .D(n22191), .CK(clk), .QN(n18254) );
  DFF_X1 avector03_reg_2__14_ ( .D(n22190), .CK(clk), .QN(n18217) );
  DFF_X1 avector03_reg_2__15_ ( .D(n22189), .CK(clk), .QN(n18180) );
  DFF_X1 avector33_reg_2__0_ ( .D(n21100), .CK(clk), .QN(n16959) );
  DFF_X1 avector33_reg_2__1_ ( .D(n21099), .CK(clk), .QN(n16922) );
  DFF_X1 avector33_reg_2__2_ ( .D(n21098), .CK(clk), .QN(n16885) );
  DFF_X1 avector33_reg_2__3_ ( .D(n21097), .CK(clk), .QN(n16848) );
  DFF_X1 avector33_reg_2__4_ ( .D(n21096), .CK(clk), .QN(n16811) );
  DFF_X1 avector33_reg_2__5_ ( .D(n21095), .CK(clk), .QN(n16774) );
  DFF_X1 avector33_reg_2__6_ ( .D(n21094), .CK(clk), .QN(n16737) );
  DFF_X1 avector33_reg_2__7_ ( .D(n21093), .CK(clk), .QN(n16700) );
  DFF_X1 avector33_reg_2__8_ ( .D(n21092), .CK(clk), .QN(n16663) );
  DFF_X1 avector33_reg_2__9_ ( .D(n21091), .CK(clk), .QN(n16626) );
  DFF_X1 avector33_reg_2__10_ ( .D(n21090), .CK(clk), .QN(n16589) );
  DFF_X1 avector33_reg_2__11_ ( .D(n21089), .CK(clk), .QN(n16552) );
  DFF_X1 avector33_reg_2__12_ ( .D(n21088), .CK(clk), .QN(n16515) );
  DFF_X1 avector33_reg_2__13_ ( .D(n21087), .CK(clk), .QN(n16478) );
  DFF_X1 avector33_reg_2__14_ ( .D(n21086), .CK(clk), .QN(n16441) );
  DFF_X1 avector33_reg_2__15_ ( .D(n21085), .CK(clk), .QN(n16404) );
  DFF_X1 avector22_reg_2__0_ ( .D(n22140), .CK(clk), .QN(n17524) );
  DFF_X1 avector22_reg_2__1_ ( .D(n22139), .CK(clk), .QN(n17487) );
  DFF_X1 avector22_reg_2__2_ ( .D(n22138), .CK(clk), .QN(n17450) );
  DFF_X1 avector22_reg_2__3_ ( .D(n22137), .CK(clk), .QN(n17413) );
  DFF_X1 avector22_reg_2__4_ ( .D(n22136), .CK(clk), .QN(n17376) );
  DFF_X1 avector22_reg_2__5_ ( .D(n22135), .CK(clk), .QN(n17339) );
  DFF_X1 avector22_reg_2__6_ ( .D(n22134), .CK(clk), .QN(n17302) );
  DFF_X1 avector22_reg_2__7_ ( .D(n22133), .CK(clk), .QN(n17265) );
  DFF_X1 avector22_reg_2__8_ ( .D(n22132), .CK(clk), .QN(n17228) );
  DFF_X1 avector22_reg_2__9_ ( .D(n22131), .CK(clk), .QN(n17191) );
  DFF_X1 avector22_reg_2__10_ ( .D(n22130), .CK(clk), .QN(n17154) );
  DFF_X1 avector22_reg_2__11_ ( .D(n22129), .CK(clk), .QN(n17117) );
  DFF_X1 avector22_reg_2__12_ ( .D(n22128), .CK(clk), .QN(n17080) );
  DFF_X1 avector22_reg_2__13_ ( .D(n22127), .CK(clk), .QN(n17043) );
  DFF_X1 avector22_reg_2__14_ ( .D(n22126), .CK(clk), .QN(n17006) );
  DFF_X1 avector22_reg_2__15_ ( .D(n22125), .CK(clk), .QN(n16969) );
  DFF_X1 avector12_reg_2__0_ ( .D(n22076), .CK(clk), .QN(n18116) );
  DFF_X1 avector12_reg_2__1_ ( .D(n22075), .CK(clk), .QN(n18079) );
  DFF_X1 avector12_reg_2__2_ ( .D(n22074), .CK(clk), .QN(n18042) );
  DFF_X1 avector12_reg_2__3_ ( .D(n22073), .CK(clk), .QN(n18005) );
  DFF_X1 avector12_reg_2__4_ ( .D(n22072), .CK(clk), .QN(n17968) );
  DFF_X1 avector12_reg_2__5_ ( .D(n22071), .CK(clk), .QN(n17931) );
  DFF_X1 avector12_reg_2__6_ ( .D(n22070), .CK(clk), .QN(n17894) );
  DFF_X1 avector12_reg_2__7_ ( .D(n22069), .CK(clk), .QN(n17857) );
  DFF_X1 avector12_reg_2__8_ ( .D(n22068), .CK(clk), .QN(n17820) );
  DFF_X1 avector12_reg_2__9_ ( .D(n22067), .CK(clk), .QN(n17783) );
  DFF_X1 avector12_reg_2__10_ ( .D(n22066), .CK(clk), .QN(n17746) );
  DFF_X1 avector12_reg_2__11_ ( .D(n22065), .CK(clk), .QN(n17709) );
  DFF_X1 avector12_reg_2__12_ ( .D(n22064), .CK(clk), .QN(n17672) );
  DFF_X1 avector12_reg_2__13_ ( .D(n22063), .CK(clk), .QN(n17635) );
  DFF_X1 avector12_reg_2__14_ ( .D(n22062), .CK(clk), .QN(n17598) );
  DFF_X1 avector12_reg_2__15_ ( .D(n22061), .CK(clk), .QN(n17561) );
  DFF_X1 avector02_reg_2__0_ ( .D(n22012), .CK(clk), .QN(n18708) );
  DFF_X1 avector02_reg_2__1_ ( .D(n22011), .CK(clk), .QN(n18671) );
  DFF_X1 avector02_reg_2__2_ ( .D(n22010), .CK(clk), .QN(n18634) );
  DFF_X1 avector02_reg_2__3_ ( .D(n22009), .CK(clk), .QN(n18597) );
  DFF_X1 avector02_reg_2__4_ ( .D(n22008), .CK(clk), .QN(n18560) );
  DFF_X1 avector02_reg_2__5_ ( .D(n22007), .CK(clk), .QN(n18523) );
  DFF_X1 avector02_reg_2__6_ ( .D(n22006), .CK(clk), .QN(n18486) );
  DFF_X1 avector02_reg_2__7_ ( .D(n22005), .CK(clk), .QN(n18449) );
  DFF_X1 avector02_reg_2__8_ ( .D(n22004), .CK(clk), .QN(n18412) );
  DFF_X1 avector02_reg_2__9_ ( .D(n22003), .CK(clk), .QN(n18375) );
  DFF_X1 avector02_reg_2__10_ ( .D(n22002), .CK(clk), .QN(n18338) );
  DFF_X1 avector02_reg_2__11_ ( .D(n22001), .CK(clk), .QN(n18301) );
  DFF_X1 avector02_reg_2__12_ ( .D(n22000), .CK(clk), .QN(n18264) );
  DFF_X1 avector02_reg_2__13_ ( .D(n21999), .CK(clk), .QN(n18227) );
  DFF_X1 avector02_reg_2__14_ ( .D(n21998), .CK(clk), .QN(n18190) );
  DFF_X1 avector02_reg_2__15_ ( .D(n21997), .CK(clk), .QN(n18153) );
  DFF_X1 avector32_reg_2__0_ ( .D(n21948), .CK(clk), .QN(n16932) );
  DFF_X1 avector32_reg_2__1_ ( .D(n21947), .CK(clk), .QN(n16895) );
  DFF_X1 avector32_reg_2__2_ ( .D(n21946), .CK(clk), .QN(n16858) );
  DFF_X1 avector32_reg_2__3_ ( .D(n21945), .CK(clk), .QN(n16821) );
  DFF_X1 avector32_reg_2__4_ ( .D(n21944), .CK(clk), .QN(n16784) );
  DFF_X1 avector32_reg_2__5_ ( .D(n21943), .CK(clk), .QN(n16747) );
  DFF_X1 avector32_reg_2__6_ ( .D(n21942), .CK(clk), .QN(n16710) );
  DFF_X1 avector32_reg_2__7_ ( .D(n21941), .CK(clk), .QN(n16673) );
  DFF_X1 avector32_reg_2__8_ ( .D(n21940), .CK(clk), .QN(n16636) );
  DFF_X1 avector32_reg_2__9_ ( .D(n21939), .CK(clk), .QN(n16599) );
  DFF_X1 avector32_reg_2__10_ ( .D(n21938), .CK(clk), .QN(n16562) );
  DFF_X1 avector32_reg_2__11_ ( .D(n21937), .CK(clk), .QN(n16525) );
  DFF_X1 avector32_reg_2__12_ ( .D(n21936), .CK(clk), .QN(n16488) );
  DFF_X1 avector32_reg_2__13_ ( .D(n21935), .CK(clk), .QN(n16451) );
  DFF_X1 avector32_reg_2__14_ ( .D(n21934), .CK(clk), .QN(n16414) );
  DFF_X1 avector32_reg_2__15_ ( .D(n21933), .CK(clk), .QN(n16377) );
  DFF_X1 avector21_reg_2__0_ ( .D(n21884), .CK(clk), .Q(n25471), .QN(n17533)
         );
  DFF_X1 avector21_reg_2__1_ ( .D(n21883), .CK(clk), .Q(n25468), .QN(n17496)
         );
  DFF_X1 avector21_reg_2__2_ ( .D(n21882), .CK(clk), .Q(n25465), .QN(n17459)
         );
  DFF_X1 avector21_reg_2__3_ ( .D(n21881), .CK(clk), .Q(n25462), .QN(n17422)
         );
  DFF_X1 avector21_reg_2__4_ ( .D(n21880), .CK(clk), .Q(n25459), .QN(n17385)
         );
  DFF_X1 avector21_reg_2__5_ ( .D(n21879), .CK(clk), .Q(n25456), .QN(n17348)
         );
  DFF_X1 avector21_reg_2__6_ ( .D(n21878), .CK(clk), .Q(n25453), .QN(n17311)
         );
  DFF_X1 avector21_reg_2__7_ ( .D(n21877), .CK(clk), .Q(n25450), .QN(n17274)
         );
  DFF_X1 avector21_reg_2__8_ ( .D(n21876), .CK(clk), .Q(n25447), .QN(n17237)
         );
  DFF_X1 avector21_reg_2__9_ ( .D(n21875), .CK(clk), .Q(n25444), .QN(n17200)
         );
  DFF_X1 avector21_reg_2__10_ ( .D(n21874), .CK(clk), .Q(n25441), .QN(n17163)
         );
  DFF_X1 avector21_reg_2__11_ ( .D(n21873), .CK(clk), .Q(n25438), .QN(n17126)
         );
  DFF_X1 avector21_reg_2__12_ ( .D(n21872), .CK(clk), .Q(n25150), .QN(n17089)
         );
  DFF_X1 avector21_reg_2__13_ ( .D(n21871), .CK(clk), .Q(n25147), .QN(n17052)
         );
  DFF_X1 avector21_reg_2__14_ ( .D(n21870), .CK(clk), .Q(n25144), .QN(n17015)
         );
  DFF_X1 avector21_reg_2__15_ ( .D(n21869), .CK(clk), .Q(n25141), .QN(n16978)
         );
  DFF_X1 avector11_reg_2__0_ ( .D(n21820), .CK(clk), .Q(n25511), .QN(n18125)
         );
  DFF_X1 avector11_reg_2__1_ ( .D(n21819), .CK(clk), .Q(n25508), .QN(n18088)
         );
  DFF_X1 avector11_reg_2__2_ ( .D(n21818), .CK(clk), .Q(n25505), .QN(n18051)
         );
  DFF_X1 avector11_reg_2__3_ ( .D(n21817), .CK(clk), .Q(n25502), .QN(n18014)
         );
  DFF_X1 avector11_reg_2__4_ ( .D(n21816), .CK(clk), .Q(n25499), .QN(n17977)
         );
  DFF_X1 avector11_reg_2__5_ ( .D(n21815), .CK(clk), .Q(n25496), .QN(n17940)
         );
  DFF_X1 avector11_reg_2__6_ ( .D(n21814), .CK(clk), .Q(n25493), .QN(n17903)
         );
  DFF_X1 avector11_reg_2__7_ ( .D(n21813), .CK(clk), .Q(n25490), .QN(n17866)
         );
  DFF_X1 avector11_reg_2__8_ ( .D(n21812), .CK(clk), .Q(n25487), .QN(n17829)
         );
  DFF_X1 avector11_reg_2__9_ ( .D(n21811), .CK(clk), .Q(n25484), .QN(n17792)
         );
  DFF_X1 avector11_reg_2__10_ ( .D(n21810), .CK(clk), .Q(n25481), .QN(n17755)
         );
  DFF_X1 avector11_reg_2__11_ ( .D(n21809), .CK(clk), .Q(n25478), .QN(n17718)
         );
  DFF_X1 avector11_reg_2__12_ ( .D(n21808), .CK(clk), .Q(n25174), .QN(n17681)
         );
  DFF_X1 avector11_reg_2__13_ ( .D(n21807), .CK(clk), .Q(n25171), .QN(n17644)
         );
  DFF_X1 avector11_reg_2__14_ ( .D(n21806), .CK(clk), .Q(n25168), .QN(n17607)
         );
  DFF_X1 avector11_reg_2__15_ ( .D(n21805), .CK(clk), .Q(n25165), .QN(n17570)
         );
  DFF_X1 avector01_reg_2__0_ ( .D(n21756), .CK(clk), .Q(n25551), .QN(n18717)
         );
  DFF_X1 avector01_reg_2__1_ ( .D(n21755), .CK(clk), .Q(n25548), .QN(n18680)
         );
  DFF_X1 avector01_reg_2__2_ ( .D(n21754), .CK(clk), .Q(n25545), .QN(n18643)
         );
  DFF_X1 avector01_reg_2__3_ ( .D(n21753), .CK(clk), .Q(n25542), .QN(n18606)
         );
  DFF_X1 avector01_reg_2__4_ ( .D(n21752), .CK(clk), .Q(n25539), .QN(n18569)
         );
  DFF_X1 avector01_reg_2__5_ ( .D(n21751), .CK(clk), .Q(n25536), .QN(n18532)
         );
  DFF_X1 avector01_reg_2__6_ ( .D(n21750), .CK(clk), .Q(n25533), .QN(n18495)
         );
  DFF_X1 avector01_reg_2__7_ ( .D(n21749), .CK(clk), .Q(n25530), .QN(n18458)
         );
  DFF_X1 avector01_reg_2__8_ ( .D(n21748), .CK(clk), .Q(n25527), .QN(n18421)
         );
  DFF_X1 avector01_reg_2__9_ ( .D(n21747), .CK(clk), .Q(n25524), .QN(n18384)
         );
  DFF_X1 avector01_reg_2__10_ ( .D(n21746), .CK(clk), .Q(n25521), .QN(n18347)
         );
  DFF_X1 avector01_reg_2__11_ ( .D(n21745), .CK(clk), .Q(n25518), .QN(n18310)
         );
  DFF_X1 avector01_reg_2__12_ ( .D(n21744), .CK(clk), .Q(n25198), .QN(n18273)
         );
  DFF_X1 avector01_reg_2__13_ ( .D(n21743), .CK(clk), .Q(n25195), .QN(n18236)
         );
  DFF_X1 avector01_reg_2__14_ ( .D(n21742), .CK(clk), .Q(n25192), .QN(n18199)
         );
  DFF_X1 avector01_reg_2__15_ ( .D(n21741), .CK(clk), .Q(n25189), .QN(n18162)
         );
  DFF_X1 avector31_reg_2__0_ ( .D(n21692), .CK(clk), .Q(n25431), .QN(n16941)
         );
  DFF_X1 avector31_reg_2__1_ ( .D(n21691), .CK(clk), .Q(n25428), .QN(n16904)
         );
  DFF_X1 avector31_reg_2__2_ ( .D(n21690), .CK(clk), .Q(n25424), .QN(n16867)
         );
  DFF_X1 avector31_reg_2__3_ ( .D(n21689), .CK(clk), .Q(n25421), .QN(n16830)
         );
  DFF_X1 avector31_reg_2__4_ ( .D(n21688), .CK(clk), .Q(n25418), .QN(n16793)
         );
  DFF_X1 avector31_reg_2__5_ ( .D(n21687), .CK(clk), .Q(n25415), .QN(n16756)
         );
  DFF_X1 avector31_reg_2__6_ ( .D(n21686), .CK(clk), .Q(n25134), .QN(n16719)
         );
  DFF_X1 avector31_reg_2__7_ ( .D(n21685), .CK(clk), .Q(n25131), .QN(n16682)
         );
  DFF_X1 avector31_reg_2__8_ ( .D(n21684), .CK(clk), .Q(n25128), .QN(n16645)
         );
  DFF_X1 avector31_reg_2__9_ ( .D(n21683), .CK(clk), .Q(n25125), .QN(n16608)
         );
  DFF_X1 avector31_reg_2__10_ ( .D(n21682), .CK(clk), .Q(n25122), .QN(n16571)
         );
  DFF_X1 avector31_reg_2__11_ ( .D(n21681), .CK(clk), .Q(n25119), .QN(n16534)
         );
  DFF_X1 avector31_reg_2__12_ ( .D(n21680), .CK(clk), .Q(n25116), .QN(n16497)
         );
  DFF_X1 avector31_reg_2__13_ ( .D(n21679), .CK(clk), .Q(n25113), .QN(n16460)
         );
  DFF_X1 avector31_reg_2__14_ ( .D(n21678), .CK(clk), .Q(n25110), .QN(n16423)
         );
  DFF_X1 avector31_reg_2__15_ ( .D(n21677), .CK(clk), .Q(n25107), .QN(n16386)
         );
  DFF_X1 avector20_reg_2__0_ ( .D(n21628), .CK(clk), .Q(n25004), .QN(n17542)
         );
  DFF_X1 avector20_reg_2__1_ ( .D(n21627), .CK(clk), .Q(n25002), .QN(n17505)
         );
  DFF_X1 avector20_reg_2__2_ ( .D(n21626), .CK(clk), .Q(n25000), .QN(n17468)
         );
  DFF_X1 avector20_reg_2__3_ ( .D(n21625), .CK(clk), .Q(n24998), .QN(n17431)
         );
  DFF_X1 avector20_reg_2__4_ ( .D(n21624), .CK(clk), .Q(n24996), .QN(n17394)
         );
  DFF_X1 avector20_reg_2__5_ ( .D(n21623), .CK(clk), .Q(n24994), .QN(n17357)
         );
  DFF_X1 avector20_reg_2__6_ ( .D(n21622), .CK(clk), .Q(n24992), .QN(n17320)
         );
  DFF_X1 avector20_reg_2__7_ ( .D(n21621), .CK(clk), .Q(n24990), .QN(n17283)
         );
  DFF_X1 avector20_reg_2__8_ ( .D(n21620), .CK(clk), .Q(n24988), .QN(n17246)
         );
  DFF_X1 avector20_reg_2__9_ ( .D(n21619), .CK(clk), .Q(n24986), .QN(n17209)
         );
  DFF_X1 avector20_reg_2__10_ ( .D(n21618), .CK(clk), .Q(n24984), .QN(n17172)
         );
  DFF_X1 avector20_reg_2__11_ ( .D(n21617), .CK(clk), .Q(n24982), .QN(n17135)
         );
  DFF_X1 avector20_reg_2__12_ ( .D(n21616), .CK(clk), .Q(n25637), .QN(n17098)
         );
  DFF_X1 avector20_reg_2__13_ ( .D(n21615), .CK(clk), .Q(n25634), .QN(n17061)
         );
  DFF_X1 avector20_reg_2__14_ ( .D(n21614), .CK(clk), .Q(n25631), .QN(n17024)
         );
  DFF_X1 avector20_reg_2__15_ ( .D(n21613), .CK(clk), .Q(n25628), .QN(n16987)
         );
  DFF_X1 avector10_reg_2__0_ ( .D(n21564), .CK(clk), .Q(n25028), .QN(n18134)
         );
  DFF_X1 avector10_reg_2__1_ ( .D(n21563), .CK(clk), .Q(n25026), .QN(n18097)
         );
  DFF_X1 avector10_reg_2__2_ ( .D(n21562), .CK(clk), .Q(n25024), .QN(n18060)
         );
  DFF_X1 avector10_reg_2__3_ ( .D(n21561), .CK(clk), .Q(n25022), .QN(n18023)
         );
  DFF_X1 avector10_reg_2__4_ ( .D(n21560), .CK(clk), .Q(n25020), .QN(n17986)
         );
  DFF_X1 avector10_reg_2__5_ ( .D(n21559), .CK(clk), .Q(n25018), .QN(n17949)
         );
  DFF_X1 avector10_reg_2__6_ ( .D(n21558), .CK(clk), .Q(n25016), .QN(n17912)
         );
  DFF_X1 avector10_reg_2__7_ ( .D(n21557), .CK(clk), .Q(n25014), .QN(n17875)
         );
  DFF_X1 avector10_reg_2__8_ ( .D(n21556), .CK(clk), .Q(n25012), .QN(n17838)
         );
  DFF_X1 avector10_reg_2__9_ ( .D(n21555), .CK(clk), .Q(n25010), .QN(n17801)
         );
  DFF_X1 avector10_reg_2__10_ ( .D(n21554), .CK(clk), .Q(n25008), .QN(n17764)
         );
  DFF_X1 avector10_reg_2__11_ ( .D(n21553), .CK(clk), .Q(n25006), .QN(n17727)
         );
  DFF_X1 avector10_reg_2__12_ ( .D(n21552), .CK(clk), .Q(n25661), .QN(n17690)
         );
  DFF_X1 avector10_reg_2__13_ ( .D(n21551), .CK(clk), .Q(n25658), .QN(n17653)
         );
  DFF_X1 avector10_reg_2__14_ ( .D(n21550), .CK(clk), .Q(n25655), .QN(n17616)
         );
  DFF_X1 avector10_reg_2__15_ ( .D(n21549), .CK(clk), .Q(n25652), .QN(n17579)
         );
  DFF_X1 avector00_reg_2__0_ ( .D(n21500), .CK(clk), .Q(n25052), .QN(n18726)
         );
  DFF_X1 avector00_reg_2__1_ ( .D(n21499), .CK(clk), .Q(n25050), .QN(n18689)
         );
  DFF_X1 avector00_reg_2__2_ ( .D(n21498), .CK(clk), .Q(n25048), .QN(n18652)
         );
  DFF_X1 avector00_reg_2__3_ ( .D(n21497), .CK(clk), .Q(n25046), .QN(n18615)
         );
  DFF_X1 avector00_reg_2__4_ ( .D(n21496), .CK(clk), .Q(n25044), .QN(n18578)
         );
  DFF_X1 avector00_reg_2__5_ ( .D(n21495), .CK(clk), .Q(n25042), .QN(n18541)
         );
  DFF_X1 avector00_reg_2__6_ ( .D(n21494), .CK(clk), .Q(n25040), .QN(n18504)
         );
  DFF_X1 avector00_reg_2__7_ ( .D(n21493), .CK(clk), .Q(n25038), .QN(n18467)
         );
  DFF_X1 avector00_reg_2__8_ ( .D(n21492), .CK(clk), .Q(n25036), .QN(n18430)
         );
  DFF_X1 avector00_reg_2__9_ ( .D(n21491), .CK(clk), .Q(n25034), .QN(n18393)
         );
  DFF_X1 avector00_reg_2__10_ ( .D(n21490), .CK(clk), .Q(n25032), .QN(n18356)
         );
  DFF_X1 avector00_reg_2__11_ ( .D(n21489), .CK(clk), .Q(n25030), .QN(n18319)
         );
  DFF_X1 avector00_reg_2__12_ ( .D(n21488), .CK(clk), .Q(n25685), .QN(n18282)
         );
  DFF_X1 avector00_reg_2__13_ ( .D(n21487), .CK(clk), .Q(n25682), .QN(n18245)
         );
  DFF_X1 avector00_reg_2__14_ ( .D(n21486), .CK(clk), .Q(n25679), .QN(n18208)
         );
  DFF_X1 avector00_reg_2__15_ ( .D(n21485), .CK(clk), .Q(n25676), .QN(n18171)
         );
  DFF_X1 avector30_reg_2__0_ ( .D(n21436), .CK(clk), .Q(n24980), .QN(n16950)
         );
  DFF_X1 avector30_reg_2__1_ ( .D(n21435), .CK(clk), .Q(n24978), .QN(n16913)
         );
  DFF_X1 avector30_reg_2__2_ ( .D(n21434), .CK(clk), .Q(n24975), .QN(n16876)
         );
  DFF_X1 avector30_reg_2__3_ ( .D(n21433), .CK(clk), .Q(n24973), .QN(n16839)
         );
  DFF_X1 avector30_reg_2__4_ ( .D(n21432), .CK(clk), .Q(n24971), .QN(n16802)
         );
  DFF_X1 avector30_reg_2__5_ ( .D(n21431), .CK(clk), .Q(n24969), .QN(n16765)
         );
  DFF_X1 avector30_reg_2__6_ ( .D(n21430), .CK(clk), .Q(n25621), .QN(n16728)
         );
  DFF_X1 avector30_reg_2__7_ ( .D(n21429), .CK(clk), .Q(n25618), .QN(n16691)
         );
  DFF_X1 avector30_reg_2__8_ ( .D(n21428), .CK(clk), .Q(n25615), .QN(n16654)
         );
  DFF_X1 avector30_reg_2__9_ ( .D(n21427), .CK(clk), .Q(n25612), .QN(n16617)
         );
  DFF_X1 avector30_reg_2__10_ ( .D(n21426), .CK(clk), .Q(n25609), .QN(n16580)
         );
  DFF_X1 avector30_reg_2__11_ ( .D(n21425), .CK(clk), .Q(n25606), .QN(n16543)
         );
  DFF_X1 avector30_reg_2__12_ ( .D(n21424), .CK(clk), .Q(n25603), .QN(n16506)
         );
  DFF_X1 avector30_reg_2__13_ ( .D(n21423), .CK(clk), .Q(n25600), .QN(n16469)
         );
  DFF_X1 avector30_reg_2__14_ ( .D(n21422), .CK(clk), .Q(n25597), .QN(n16432)
         );
  DFF_X1 avector30_reg_2__15_ ( .D(n21421), .CK(clk), .Q(n25594), .QN(n16395)
         );
  DFF_X1 avector23_reg_4__0_ ( .D(n22364), .CK(clk), .Q(n25469), .QN(n17556)
         );
  DFF_X1 avector23_reg_4__1_ ( .D(n22363), .CK(clk), .Q(n25466), .QN(n17519)
         );
  DFF_X1 avector23_reg_4__2_ ( .D(n22362), .CK(clk), .Q(n25463), .QN(n17482)
         );
  DFF_X1 avector23_reg_4__3_ ( .D(n22361), .CK(clk), .Q(n25460), .QN(n17445)
         );
  DFF_X1 avector23_reg_4__4_ ( .D(n22360), .CK(clk), .Q(n25457), .QN(n17408)
         );
  DFF_X1 avector23_reg_4__5_ ( .D(n22359), .CK(clk), .Q(n25454), .QN(n17371)
         );
  DFF_X1 avector23_reg_4__6_ ( .D(n22358), .CK(clk), .Q(n25451), .QN(n17334)
         );
  DFF_X1 avector23_reg_4__7_ ( .D(n22357), .CK(clk), .Q(n25448), .QN(n17297)
         );
  DFF_X1 avector23_reg_4__8_ ( .D(n22356), .CK(clk), .Q(n25445), .QN(n17260)
         );
  DFF_X1 avector23_reg_4__9_ ( .D(n22355), .CK(clk), .Q(n25442), .QN(n17223)
         );
  DFF_X1 avector23_reg_4__10_ ( .D(n22354), .CK(clk), .Q(n25439), .QN(n17186)
         );
  DFF_X1 avector23_reg_4__11_ ( .D(n22353), .CK(clk), .Q(n25436), .QN(n17149)
         );
  DFF_X1 avector23_reg_4__12_ ( .D(n22352), .CK(clk), .Q(n25435), .QN(n17112)
         );
  DFF_X1 avector23_reg_4__13_ ( .D(n22351), .CK(clk), .Q(n25434), .QN(n17075)
         );
  DFF_X1 avector23_reg_4__14_ ( .D(n22350), .CK(clk), .Q(n25433), .QN(n17038)
         );
  DFF_X1 avector23_reg_4__15_ ( .D(n22349), .CK(clk), .Q(n25432), .QN(n17001)
         );
  DFF_X1 avector13_reg_4__0_ ( .D(n22300), .CK(clk), .Q(n25509), .QN(n18148)
         );
  DFF_X1 avector13_reg_4__1_ ( .D(n22299), .CK(clk), .Q(n25506), .QN(n18111)
         );
  DFF_X1 avector13_reg_4__2_ ( .D(n22298), .CK(clk), .Q(n25503), .QN(n18074)
         );
  DFF_X1 avector13_reg_4__3_ ( .D(n22297), .CK(clk), .Q(n25500), .QN(n18037)
         );
  DFF_X1 avector13_reg_4__4_ ( .D(n22296), .CK(clk), .Q(n25497), .QN(n18000)
         );
  DFF_X1 avector13_reg_4__5_ ( .D(n22295), .CK(clk), .Q(n25494), .QN(n17963)
         );
  DFF_X1 avector13_reg_4__6_ ( .D(n22294), .CK(clk), .Q(n25491), .QN(n17926)
         );
  DFF_X1 avector13_reg_4__7_ ( .D(n22293), .CK(clk), .Q(n25488), .QN(n17889)
         );
  DFF_X1 avector13_reg_4__8_ ( .D(n22292), .CK(clk), .Q(n25485), .QN(n17852)
         );
  DFF_X1 avector13_reg_4__9_ ( .D(n22291), .CK(clk), .Q(n25482), .QN(n17815)
         );
  DFF_X1 avector13_reg_4__10_ ( .D(n22290), .CK(clk), .Q(n25479), .QN(n17778)
         );
  DFF_X1 avector13_reg_4__11_ ( .D(n22289), .CK(clk), .Q(n25476), .QN(n17741)
         );
  DFF_X1 avector13_reg_4__12_ ( .D(n22288), .CK(clk), .Q(n25475), .QN(n17704)
         );
  DFF_X1 avector13_reg_4__13_ ( .D(n22287), .CK(clk), .Q(n25474), .QN(n17667)
         );
  DFF_X1 avector13_reg_4__14_ ( .D(n22286), .CK(clk), .Q(n25473), .QN(n17630)
         );
  DFF_X1 avector13_reg_4__15_ ( .D(n22285), .CK(clk), .Q(n25472), .QN(n17593)
         );
  DFF_X1 avector03_reg_4__0_ ( .D(n22236), .CK(clk), .Q(n25549), .QN(n18740)
         );
  DFF_X1 avector03_reg_4__1_ ( .D(n22235), .CK(clk), .Q(n25546), .QN(n18703)
         );
  DFF_X1 avector03_reg_4__2_ ( .D(n22234), .CK(clk), .Q(n25543), .QN(n18666)
         );
  DFF_X1 avector03_reg_4__3_ ( .D(n22233), .CK(clk), .Q(n25540), .QN(n18629)
         );
  DFF_X1 avector03_reg_4__4_ ( .D(n22232), .CK(clk), .Q(n25537), .QN(n18592)
         );
  DFF_X1 avector03_reg_4__5_ ( .D(n22231), .CK(clk), .Q(n25534), .QN(n18555)
         );
  DFF_X1 avector03_reg_4__6_ ( .D(n22230), .CK(clk), .Q(n25531), .QN(n18518)
         );
  DFF_X1 avector03_reg_4__7_ ( .D(n22229), .CK(clk), .Q(n25528), .QN(n18481)
         );
  DFF_X1 avector03_reg_4__8_ ( .D(n22228), .CK(clk), .Q(n25525), .QN(n18444)
         );
  DFF_X1 avector03_reg_4__9_ ( .D(n22227), .CK(clk), .Q(n25522), .QN(n18407)
         );
  DFF_X1 avector03_reg_4__10_ ( .D(n22226), .CK(clk), .Q(n25519), .QN(n18370)
         );
  DFF_X1 avector03_reg_4__11_ ( .D(n22225), .CK(clk), .Q(n25516), .QN(n18333)
         );
  DFF_X1 avector03_reg_4__12_ ( .D(n22224), .CK(clk), .Q(n25515), .QN(n18296)
         );
  DFF_X1 avector03_reg_4__13_ ( .D(n22223), .CK(clk), .Q(n25514), .QN(n18259)
         );
  DFF_X1 avector03_reg_4__14_ ( .D(n22222), .CK(clk), .Q(n25513), .QN(n18222)
         );
  DFF_X1 avector03_reg_4__15_ ( .D(n22221), .CK(clk), .Q(n25512), .QN(n18185)
         );
  DFF_X1 avector33_reg_4__0_ ( .D(n21132), .CK(clk), .Q(n25429), .QN(n16964)
         );
  DFF_X1 avector33_reg_4__1_ ( .D(n21131), .CK(clk), .Q(n25426), .QN(n16927)
         );
  DFF_X1 avector33_reg_4__2_ ( .D(n21130), .CK(clk), .Q(n25422), .QN(n16890)
         );
  DFF_X1 avector33_reg_4__3_ ( .D(n21129), .CK(clk), .Q(n25419), .QN(n16853)
         );
  DFF_X1 avector33_reg_4__4_ ( .D(n21128), .CK(clk), .Q(n25416), .QN(n16816)
         );
  DFF_X1 avector33_reg_4__5_ ( .D(n21127), .CK(clk), .Q(n25413), .QN(n16779)
         );
  DFF_X1 avector33_reg_4__6_ ( .D(n21126), .CK(clk), .Q(n25411), .QN(n16742)
         );
  DFF_X1 avector33_reg_4__7_ ( .D(n21125), .CK(clk), .Q(n25410), .QN(n16705)
         );
  DFF_X1 avector33_reg_4__8_ ( .D(n21124), .CK(clk), .Q(n25409), .QN(n16668)
         );
  DFF_X1 avector33_reg_4__9_ ( .D(n21123), .CK(clk), .Q(n25408), .QN(n16631)
         );
  DFF_X1 avector33_reg_4__10_ ( .D(n21122), .CK(clk), .Q(n25407), .QN(n16594)
         );
  DFF_X1 avector33_reg_4__11_ ( .D(n21121), .CK(clk), .Q(n25406), .QN(n16557)
         );
  DFF_X1 avector33_reg_4__12_ ( .D(n21120), .CK(clk), .Q(n25405), .QN(n16520)
         );
  DFF_X1 avector33_reg_4__13_ ( .D(n21119), .CK(clk), .Q(n25404), .QN(n16483)
         );
  DFF_X1 avector33_reg_4__14_ ( .D(n21118), .CK(clk), .Q(n25403), .QN(n16446)
         );
  DFF_X1 avector33_reg_4__15_ ( .D(n21117), .CK(clk), .Q(n25402), .QN(n16409)
         );
  DFF_X1 avector22_reg_4__0_ ( .D(n22172), .CK(clk), .QN(n17529) );
  DFF_X1 avector22_reg_4__1_ ( .D(n22171), .CK(clk), .QN(n17492) );
  DFF_X1 avector22_reg_4__2_ ( .D(n22170), .CK(clk), .QN(n17455) );
  DFF_X1 avector22_reg_4__3_ ( .D(n22169), .CK(clk), .QN(n17418) );
  DFF_X1 avector22_reg_4__4_ ( .D(n22168), .CK(clk), .QN(n17381) );
  DFF_X1 avector22_reg_4__5_ ( .D(n22167), .CK(clk), .QN(n17344) );
  DFF_X1 avector22_reg_4__6_ ( .D(n22166), .CK(clk), .QN(n17307) );
  DFF_X1 avector22_reg_4__7_ ( .D(n22165), .CK(clk), .QN(n17270) );
  DFF_X1 avector22_reg_4__8_ ( .D(n22164), .CK(clk), .QN(n17233) );
  DFF_X1 avector22_reg_4__9_ ( .D(n22163), .CK(clk), .QN(n17196) );
  DFF_X1 avector22_reg_4__10_ ( .D(n22162), .CK(clk), .QN(n17159) );
  DFF_X1 avector22_reg_4__11_ ( .D(n22161), .CK(clk), .QN(n17122) );
  DFF_X1 avector22_reg_4__12_ ( .D(n22160), .CK(clk), .QN(n17085) );
  DFF_X1 avector22_reg_4__13_ ( .D(n22159), .CK(clk), .QN(n17048) );
  DFF_X1 avector22_reg_4__14_ ( .D(n22158), .CK(clk), .QN(n17011) );
  DFF_X1 avector22_reg_4__15_ ( .D(n22157), .CK(clk), .QN(n16974) );
  DFF_X1 avector12_reg_4__0_ ( .D(n22108), .CK(clk), .QN(n18121) );
  DFF_X1 avector12_reg_4__1_ ( .D(n22107), .CK(clk), .QN(n18084) );
  DFF_X1 avector12_reg_4__2_ ( .D(n22106), .CK(clk), .QN(n18047) );
  DFF_X1 avector12_reg_4__3_ ( .D(n22105), .CK(clk), .QN(n18010) );
  DFF_X1 avector12_reg_4__4_ ( .D(n22104), .CK(clk), .QN(n17973) );
  DFF_X1 avector12_reg_4__5_ ( .D(n22103), .CK(clk), .QN(n17936) );
  DFF_X1 avector12_reg_4__6_ ( .D(n22102), .CK(clk), .QN(n17899) );
  DFF_X1 avector12_reg_4__7_ ( .D(n22101), .CK(clk), .QN(n17862) );
  DFF_X1 avector12_reg_4__8_ ( .D(n22100), .CK(clk), .QN(n17825) );
  DFF_X1 avector12_reg_4__9_ ( .D(n22099), .CK(clk), .QN(n17788) );
  DFF_X1 avector12_reg_4__10_ ( .D(n22098), .CK(clk), .QN(n17751) );
  DFF_X1 avector12_reg_4__11_ ( .D(n22097), .CK(clk), .QN(n17714) );
  DFF_X1 avector12_reg_4__12_ ( .D(n22096), .CK(clk), .QN(n17677) );
  DFF_X1 avector12_reg_4__13_ ( .D(n22095), .CK(clk), .QN(n17640) );
  DFF_X1 avector12_reg_4__14_ ( .D(n22094), .CK(clk), .QN(n17603) );
  DFF_X1 avector12_reg_4__15_ ( .D(n22093), .CK(clk), .QN(n17566) );
  DFF_X1 avector02_reg_4__0_ ( .D(n22044), .CK(clk), .QN(n18713) );
  DFF_X1 avector02_reg_4__1_ ( .D(n22043), .CK(clk), .QN(n18676) );
  DFF_X1 avector02_reg_4__2_ ( .D(n22042), .CK(clk), .QN(n18639) );
  DFF_X1 avector02_reg_4__3_ ( .D(n22041), .CK(clk), .QN(n18602) );
  DFF_X1 avector02_reg_4__4_ ( .D(n22040), .CK(clk), .QN(n18565) );
  DFF_X1 avector02_reg_4__5_ ( .D(n22039), .CK(clk), .QN(n18528) );
  DFF_X1 avector02_reg_4__6_ ( .D(n22038), .CK(clk), .QN(n18491) );
  DFF_X1 avector02_reg_4__7_ ( .D(n22037), .CK(clk), .QN(n18454) );
  DFF_X1 avector02_reg_4__8_ ( .D(n22036), .CK(clk), .QN(n18417) );
  DFF_X1 avector02_reg_4__9_ ( .D(n22035), .CK(clk), .QN(n18380) );
  DFF_X1 avector02_reg_4__10_ ( .D(n22034), .CK(clk), .QN(n18343) );
  DFF_X1 avector02_reg_4__11_ ( .D(n22033), .CK(clk), .QN(n18306) );
  DFF_X1 avector02_reg_4__12_ ( .D(n22032), .CK(clk), .QN(n18269) );
  DFF_X1 avector02_reg_4__13_ ( .D(n22031), .CK(clk), .QN(n18232) );
  DFF_X1 avector02_reg_4__14_ ( .D(n22030), .CK(clk), .QN(n18195) );
  DFF_X1 avector02_reg_4__15_ ( .D(n22029), .CK(clk), .QN(n18158) );
  DFF_X1 avector32_reg_4__0_ ( .D(n21980), .CK(clk), .QN(n16937) );
  DFF_X1 avector32_reg_4__1_ ( .D(n21979), .CK(clk), .QN(n16900) );
  DFF_X1 avector32_reg_4__2_ ( .D(n21978), .CK(clk), .QN(n16863) );
  DFF_X1 avector32_reg_4__3_ ( .D(n21977), .CK(clk), .QN(n16826) );
  DFF_X1 avector32_reg_4__4_ ( .D(n21976), .CK(clk), .QN(n16789) );
  DFF_X1 avector32_reg_4__5_ ( .D(n21975), .CK(clk), .QN(n16752) );
  DFF_X1 avector32_reg_4__6_ ( .D(n21974), .CK(clk), .QN(n16715) );
  DFF_X1 avector32_reg_4__7_ ( .D(n21973), .CK(clk), .QN(n16678) );
  DFF_X1 avector32_reg_4__8_ ( .D(n21972), .CK(clk), .QN(n16641) );
  DFF_X1 avector32_reg_4__9_ ( .D(n21971), .CK(clk), .QN(n16604) );
  DFF_X1 avector32_reg_4__10_ ( .D(n21970), .CK(clk), .QN(n16567) );
  DFF_X1 avector32_reg_4__11_ ( .D(n21969), .CK(clk), .QN(n16530) );
  DFF_X1 avector32_reg_4__12_ ( .D(n21968), .CK(clk), .QN(n16493) );
  DFF_X1 avector32_reg_4__13_ ( .D(n21967), .CK(clk), .QN(n16456) );
  DFF_X1 avector32_reg_4__14_ ( .D(n21966), .CK(clk), .QN(n16419) );
  DFF_X1 avector32_reg_4__15_ ( .D(n21965), .CK(clk), .QN(n16382) );
  DFF_X1 avector21_reg_4__0_ ( .D(n21916), .CK(clk), .Q(n25162), .QN(n17538)
         );
  DFF_X1 avector21_reg_4__1_ ( .D(n21915), .CK(clk), .Q(n25161), .QN(n17501)
         );
  DFF_X1 avector21_reg_4__2_ ( .D(n21914), .CK(clk), .Q(n25160), .QN(n17464)
         );
  DFF_X1 avector21_reg_4__3_ ( .D(n21913), .CK(clk), .Q(n25159), .QN(n17427)
         );
  DFF_X1 avector21_reg_4__4_ ( .D(n21912), .CK(clk), .Q(n25158), .QN(n17390)
         );
  DFF_X1 avector21_reg_4__5_ ( .D(n21911), .CK(clk), .Q(n25157), .QN(n17353)
         );
  DFF_X1 avector21_reg_4__6_ ( .D(n21910), .CK(clk), .Q(n25156), .QN(n17316)
         );
  DFF_X1 avector21_reg_4__7_ ( .D(n21909), .CK(clk), .Q(n25155), .QN(n17279)
         );
  DFF_X1 avector21_reg_4__8_ ( .D(n21908), .CK(clk), .Q(n25154), .QN(n17242)
         );
  DFF_X1 avector21_reg_4__9_ ( .D(n21907), .CK(clk), .Q(n25153), .QN(n17205)
         );
  DFF_X1 avector21_reg_4__10_ ( .D(n21906), .CK(clk), .Q(n25152), .QN(n17168)
         );
  DFF_X1 avector21_reg_4__11_ ( .D(n21905), .CK(clk), .Q(n25151), .QN(n17131)
         );
  DFF_X1 avector21_reg_4__12_ ( .D(n21904), .CK(clk), .Q(n25148), .QN(n17094)
         );
  DFF_X1 avector21_reg_4__13_ ( .D(n21903), .CK(clk), .Q(n25145), .QN(n17057)
         );
  DFF_X1 avector21_reg_4__14_ ( .D(n21902), .CK(clk), .Q(n25142), .QN(n17020)
         );
  DFF_X1 avector21_reg_4__15_ ( .D(n21901), .CK(clk), .Q(n25139), .QN(n16983)
         );
  DFF_X1 avector11_reg_4__0_ ( .D(n21852), .CK(clk), .Q(n25186), .QN(n18130)
         );
  DFF_X1 avector11_reg_4__1_ ( .D(n21851), .CK(clk), .Q(n25185), .QN(n18093)
         );
  DFF_X1 avector11_reg_4__2_ ( .D(n21850), .CK(clk), .Q(n25184), .QN(n18056)
         );
  DFF_X1 avector11_reg_4__3_ ( .D(n21849), .CK(clk), .Q(n25183), .QN(n18019)
         );
  DFF_X1 avector11_reg_4__4_ ( .D(n21848), .CK(clk), .Q(n25182), .QN(n17982)
         );
  DFF_X1 avector11_reg_4__5_ ( .D(n21847), .CK(clk), .Q(n25181), .QN(n17945)
         );
  DFF_X1 avector11_reg_4__6_ ( .D(n21846), .CK(clk), .Q(n25180), .QN(n17908)
         );
  DFF_X1 avector11_reg_4__7_ ( .D(n21845), .CK(clk), .Q(n25179), .QN(n17871)
         );
  DFF_X1 avector11_reg_4__8_ ( .D(n21844), .CK(clk), .Q(n25178), .QN(n17834)
         );
  DFF_X1 avector11_reg_4__9_ ( .D(n21843), .CK(clk), .Q(n25177), .QN(n17797)
         );
  DFF_X1 avector11_reg_4__10_ ( .D(n21842), .CK(clk), .Q(n25176), .QN(n17760)
         );
  DFF_X1 avector11_reg_4__11_ ( .D(n21841), .CK(clk), .Q(n25175), .QN(n17723)
         );
  DFF_X1 avector11_reg_4__12_ ( .D(n21840), .CK(clk), .Q(n25172), .QN(n17686)
         );
  DFF_X1 avector11_reg_4__13_ ( .D(n21839), .CK(clk), .Q(n25169), .QN(n17649)
         );
  DFF_X1 avector11_reg_4__14_ ( .D(n21838), .CK(clk), .Q(n25166), .QN(n17612)
         );
  DFF_X1 avector11_reg_4__15_ ( .D(n21837), .CK(clk), .Q(n25163), .QN(n17575)
         );
  DFF_X1 avector01_reg_4__0_ ( .D(n21788), .CK(clk), .Q(n25210), .QN(n18722)
         );
  DFF_X1 avector01_reg_4__1_ ( .D(n21787), .CK(clk), .Q(n25209), .QN(n18685)
         );
  DFF_X1 avector01_reg_4__2_ ( .D(n21786), .CK(clk), .Q(n25208), .QN(n18648)
         );
  DFF_X1 avector01_reg_4__3_ ( .D(n21785), .CK(clk), .Q(n25207), .QN(n18611)
         );
  DFF_X1 avector01_reg_4__4_ ( .D(n21784), .CK(clk), .Q(n25206), .QN(n18574)
         );
  DFF_X1 avector01_reg_4__5_ ( .D(n21783), .CK(clk), .Q(n25205), .QN(n18537)
         );
  DFF_X1 avector01_reg_4__6_ ( .D(n21782), .CK(clk), .Q(n25204), .QN(n18500)
         );
  DFF_X1 avector01_reg_4__7_ ( .D(n21781), .CK(clk), .Q(n25203), .QN(n18463)
         );
  DFF_X1 avector01_reg_4__8_ ( .D(n21780), .CK(clk), .Q(n25202), .QN(n18426)
         );
  DFF_X1 avector01_reg_4__9_ ( .D(n21779), .CK(clk), .Q(n25201), .QN(n18389)
         );
  DFF_X1 avector01_reg_4__10_ ( .D(n21778), .CK(clk), .Q(n25200), .QN(n18352)
         );
  DFF_X1 avector01_reg_4__11_ ( .D(n21777), .CK(clk), .Q(n25199), .QN(n18315)
         );
  DFF_X1 avector01_reg_4__12_ ( .D(n21776), .CK(clk), .Q(n25196), .QN(n18278)
         );
  DFF_X1 avector01_reg_4__13_ ( .D(n21775), .CK(clk), .Q(n25193), .QN(n18241)
         );
  DFF_X1 avector01_reg_4__14_ ( .D(n21774), .CK(clk), .Q(n25190), .QN(n18204)
         );
  DFF_X1 avector01_reg_4__15_ ( .D(n21773), .CK(clk), .Q(n25187), .QN(n18167)
         );
  DFF_X1 avector31_reg_4__0_ ( .D(n21724), .CK(clk), .Q(n25138), .QN(n16946)
         );
  DFF_X1 avector31_reg_4__1_ ( .D(n21723), .CK(clk), .Q(n25425), .QN(n16909)
         );
  DFF_X1 avector31_reg_4__2_ ( .D(n21722), .CK(clk), .Q(n25137), .QN(n16872)
         );
  DFF_X1 avector31_reg_4__3_ ( .D(n21721), .CK(clk), .Q(n25136), .QN(n16835)
         );
  DFF_X1 avector31_reg_4__4_ ( .D(n21720), .CK(clk), .Q(n25135), .QN(n16798)
         );
  DFF_X1 avector31_reg_4__5_ ( .D(n21719), .CK(clk), .Q(n25412), .QN(n16761)
         );
  DFF_X1 avector31_reg_4__6_ ( .D(n21718), .CK(clk), .Q(n25132), .QN(n16724)
         );
  DFF_X1 avector31_reg_4__7_ ( .D(n21717), .CK(clk), .Q(n25129), .QN(n16687)
         );
  DFF_X1 avector31_reg_4__8_ ( .D(n21716), .CK(clk), .Q(n25126), .QN(n16650)
         );
  DFF_X1 avector31_reg_4__9_ ( .D(n21715), .CK(clk), .Q(n25123), .QN(n16613)
         );
  DFF_X1 avector31_reg_4__10_ ( .D(n21714), .CK(clk), .Q(n25120), .QN(n16576)
         );
  DFF_X1 avector31_reg_4__11_ ( .D(n21713), .CK(clk), .Q(n25117), .QN(n16539)
         );
  DFF_X1 avector31_reg_4__12_ ( .D(n21712), .CK(clk), .Q(n25114), .QN(n16502)
         );
  DFF_X1 avector31_reg_4__13_ ( .D(n21711), .CK(clk), .Q(n25111), .QN(n16465)
         );
  DFF_X1 avector31_reg_4__14_ ( .D(n21710), .CK(clk), .Q(n25108), .QN(n16428)
         );
  DFF_X1 avector31_reg_4__15_ ( .D(n21709), .CK(clk), .Q(n25105), .QN(n16391)
         );
  DFF_X1 avector20_reg_4__0_ ( .D(n21660), .CK(clk), .Q(n25649), .QN(n17547)
         );
  DFF_X1 avector20_reg_4__1_ ( .D(n21659), .CK(clk), .Q(n25648), .QN(n17510)
         );
  DFF_X1 avector20_reg_4__2_ ( .D(n21658), .CK(clk), .Q(n25647), .QN(n17473)
         );
  DFF_X1 avector20_reg_4__3_ ( .D(n21657), .CK(clk), .Q(n25646), .QN(n17436)
         );
  DFF_X1 avector20_reg_4__4_ ( .D(n21656), .CK(clk), .Q(n25645), .QN(n17399)
         );
  DFF_X1 avector20_reg_4__5_ ( .D(n21655), .CK(clk), .Q(n25644), .QN(n17362)
         );
  DFF_X1 avector20_reg_4__6_ ( .D(n21654), .CK(clk), .Q(n25643), .QN(n17325)
         );
  DFF_X1 avector20_reg_4__7_ ( .D(n21653), .CK(clk), .Q(n25642), .QN(n17288)
         );
  DFF_X1 avector20_reg_4__8_ ( .D(n21652), .CK(clk), .Q(n25641), .QN(n17251)
         );
  DFF_X1 avector20_reg_4__9_ ( .D(n21651), .CK(clk), .Q(n25640), .QN(n17214)
         );
  DFF_X1 avector20_reg_4__10_ ( .D(n21650), .CK(clk), .Q(n25639), .QN(n17177)
         );
  DFF_X1 avector20_reg_4__11_ ( .D(n21649), .CK(clk), .Q(n25638), .QN(n17140)
         );
  DFF_X1 avector20_reg_4__12_ ( .D(n21648), .CK(clk), .Q(n25635), .QN(n17103)
         );
  DFF_X1 avector20_reg_4__13_ ( .D(n21647), .CK(clk), .Q(n25632), .QN(n17066)
         );
  DFF_X1 avector20_reg_4__14_ ( .D(n21646), .CK(clk), .Q(n25629), .QN(n17029)
         );
  DFF_X1 avector20_reg_4__15_ ( .D(n21645), .CK(clk), .Q(n25626), .QN(n16992)
         );
  DFF_X1 avector10_reg_4__0_ ( .D(n21596), .CK(clk), .Q(n25673), .QN(n18139)
         );
  DFF_X1 avector10_reg_4__1_ ( .D(n21595), .CK(clk), .Q(n25672), .QN(n18102)
         );
  DFF_X1 avector10_reg_4__2_ ( .D(n21594), .CK(clk), .Q(n25671), .QN(n18065)
         );
  DFF_X1 avector10_reg_4__3_ ( .D(n21593), .CK(clk), .Q(n25670), .QN(n18028)
         );
  DFF_X1 avector10_reg_4__4_ ( .D(n21592), .CK(clk), .Q(n25669), .QN(n17991)
         );
  DFF_X1 avector10_reg_4__5_ ( .D(n21591), .CK(clk), .Q(n25668), .QN(n17954)
         );
  DFF_X1 avector10_reg_4__6_ ( .D(n21590), .CK(clk), .Q(n25667), .QN(n17917)
         );
  DFF_X1 avector10_reg_4__7_ ( .D(n21589), .CK(clk), .Q(n25666), .QN(n17880)
         );
  DFF_X1 avector10_reg_4__8_ ( .D(n21588), .CK(clk), .Q(n25665), .QN(n17843)
         );
  DFF_X1 avector10_reg_4__9_ ( .D(n21587), .CK(clk), .Q(n25664), .QN(n17806)
         );
  DFF_X1 avector10_reg_4__10_ ( .D(n21586), .CK(clk), .Q(n25663), .QN(n17769)
         );
  DFF_X1 avector10_reg_4__11_ ( .D(n21585), .CK(clk), .Q(n25662), .QN(n17732)
         );
  DFF_X1 avector10_reg_4__12_ ( .D(n21584), .CK(clk), .Q(n25659), .QN(n17695)
         );
  DFF_X1 avector10_reg_4__13_ ( .D(n21583), .CK(clk), .Q(n25656), .QN(n17658)
         );
  DFF_X1 avector10_reg_4__14_ ( .D(n21582), .CK(clk), .Q(n25653), .QN(n17621)
         );
  DFF_X1 avector10_reg_4__15_ ( .D(n21581), .CK(clk), .Q(n25650), .QN(n17584)
         );
  DFF_X1 avector00_reg_4__0_ ( .D(n21532), .CK(clk), .Q(n25697), .QN(n18731)
         );
  DFF_X1 avector00_reg_4__1_ ( .D(n21531), .CK(clk), .Q(n25696), .QN(n18694)
         );
  DFF_X1 avector00_reg_4__2_ ( .D(n21530), .CK(clk), .Q(n25695), .QN(n18657)
         );
  DFF_X1 avector00_reg_4__3_ ( .D(n21529), .CK(clk), .Q(n25694), .QN(n18620)
         );
  DFF_X1 avector00_reg_4__4_ ( .D(n21528), .CK(clk), .Q(n25693), .QN(n18583)
         );
  DFF_X1 avector00_reg_4__5_ ( .D(n21527), .CK(clk), .Q(n25692), .QN(n18546)
         );
  DFF_X1 avector00_reg_4__6_ ( .D(n21526), .CK(clk), .Q(n25691), .QN(n18509)
         );
  DFF_X1 avector00_reg_4__7_ ( .D(n21525), .CK(clk), .Q(n25690), .QN(n18472)
         );
  DFF_X1 avector00_reg_4__8_ ( .D(n21524), .CK(clk), .Q(n25689), .QN(n18435)
         );
  DFF_X1 avector00_reg_4__9_ ( .D(n21523), .CK(clk), .Q(n25688), .QN(n18398)
         );
  DFF_X1 avector00_reg_4__10_ ( .D(n21522), .CK(clk), .Q(n25687), .QN(n18361)
         );
  DFF_X1 avector00_reg_4__11_ ( .D(n21521), .CK(clk), .Q(n25686), .QN(n18324)
         );
  DFF_X1 avector00_reg_4__12_ ( .D(n21520), .CK(clk), .Q(n25683), .QN(n18287)
         );
  DFF_X1 avector00_reg_4__13_ ( .D(n21519), .CK(clk), .Q(n25680), .QN(n18250)
         );
  DFF_X1 avector00_reg_4__14_ ( .D(n21518), .CK(clk), .Q(n25677), .QN(n18213)
         );
  DFF_X1 avector00_reg_4__15_ ( .D(n21517), .CK(clk), .Q(n25674), .QN(n18176)
         );
  DFF_X1 avector30_reg_4__0_ ( .D(n21468), .CK(clk), .Q(n25625), .QN(n16955)
         );
  DFF_X1 avector30_reg_4__1_ ( .D(n21467), .CK(clk), .Q(n24976), .QN(n16918)
         );
  DFF_X1 avector30_reg_4__2_ ( .D(n21466), .CK(clk), .Q(n25624), .QN(n16881)
         );
  DFF_X1 avector30_reg_4__3_ ( .D(n21465), .CK(clk), .Q(n25623), .QN(n16844)
         );
  DFF_X1 avector30_reg_4__4_ ( .D(n21464), .CK(clk), .Q(n25622), .QN(n16807)
         );
  DFF_X1 avector30_reg_4__5_ ( .D(n21463), .CK(clk), .Q(n24967), .QN(n16770)
         );
  DFF_X1 avector30_reg_4__6_ ( .D(n21462), .CK(clk), .Q(n25619), .QN(n16733)
         );
  DFF_X1 avector30_reg_4__7_ ( .D(n21461), .CK(clk), .Q(n25616), .QN(n16696)
         );
  DFF_X1 avector30_reg_4__8_ ( .D(n21460), .CK(clk), .Q(n25613), .QN(n16659)
         );
  DFF_X1 avector30_reg_4__9_ ( .D(n21459), .CK(clk), .Q(n25610), .QN(n16622)
         );
  DFF_X1 avector30_reg_4__10_ ( .D(n21458), .CK(clk), .Q(n25607), .QN(n16585)
         );
  DFF_X1 avector30_reg_4__11_ ( .D(n21457), .CK(clk), .Q(n25604), .QN(n16548)
         );
  DFF_X1 avector30_reg_4__12_ ( .D(n21456), .CK(clk), .Q(n25601), .QN(n16511)
         );
  DFF_X1 avector30_reg_4__13_ ( .D(n21455), .CK(clk), .Q(n25598), .QN(n16474)
         );
  DFF_X1 avector30_reg_4__14_ ( .D(n21454), .CK(clk), .Q(n25595), .QN(n16437)
         );
  DFF_X1 avector30_reg_4__15_ ( .D(n21453), .CK(clk), .Q(n25592), .QN(n16400)
         );
  DFF_X1 select_reg_0_ ( .D(n23519), .CK(clk), .Q(n24890), .QN(n22398) );
  DFF_X1 select_reg_1_ ( .D(n23518), .CK(clk), .Q(n25245), .QN(n22397) );
  DFF_X1 select_reg_2_ ( .D(n23517), .CK(clk), .QN(n22396) );
  DFF_X1 select_reg_3_ ( .D(n23516), .CK(clk), .Q(n25246), .QN(n22395) );
  DFF_X1 bitselect2_reg_0_ ( .D(n23450), .CK(clk), .QN(n22406) );
  DFF_X1 zcount_reg_0_ ( .D(n23446), .CK(clk), .Q(n25253), .QN(n22403) );
  DFF_X1 zcount_reg_1_ ( .D(n21084), .CK(clk), .Q(n24887), .QN(n22402) );
  DFF_X1 zcount_reg_2_ ( .D(n23445), .CK(clk), .Q(n24896), .QN(n22401) );
  DFF_X1 zcount_reg_3_ ( .D(n23444), .CK(clk), .Q(n25257), .QN(n22400) );
  DFF_X1 bitselect2_reg_1_ ( .D(n23449), .CK(clk), .Q(n25104), .QN(n22405) );
  DFF_X1 bitselect2_reg_2_ ( .D(n23448), .CK(clk), .Q(n25401), .QN(n22404) );
  DFF_X1 m_reg_15_ ( .D(n20571), .CK(clk), .Q(n5056), .QN(n20539) );
  DFF_X1 m_reg_14_ ( .D(n20570), .CK(clk), .Q(n5055), .QN(n20538) );
  DFF_X1 m_reg_13_ ( .D(n20569), .CK(clk), .Q(n5054), .QN(n20537) );
  DFF_X1 m_reg_12_ ( .D(n20568), .CK(clk), .Q(n5053), .QN(n20536) );
  DFF_X1 m_reg_11_ ( .D(n20567), .CK(clk), .Q(n5052), .QN(n20535) );
  DFF_X1 m_reg_10_ ( .D(n20566), .CK(clk), .Q(n5051), .QN(n20534) );
  DFF_X1 m_reg_9_ ( .D(n20565), .CK(clk), .Q(n5050), .QN(n20533) );
  DFF_X1 m_reg_8_ ( .D(n20564), .CK(clk), .Q(n5049), .QN(n20532) );
  DFF_X1 m_reg_0_ ( .D(n20556), .CK(clk), .Q(n5041), .QN(n20524) );
  DFF_X1 count_out_reg_1_ ( .D(n23432), .CK(clk), .Q(n24894), .QN(n22421) );
  DFF_X1 count_out_reg_2_ ( .D(n23431), .CK(clk), .Q(n25255), .QN(n22420) );
  DFF_X1 bvector3_reg_5__0_ ( .D(n21418), .CK(clk), .QN(n18791) );
  DFF_X1 bvector3_reg_5__1_ ( .D(n21417), .CK(clk), .QN(n18828) );
  DFF_X1 bvector3_reg_5__2_ ( .D(n21416), .CK(clk), .QN(n18865) );
  DFF_X1 bvector3_reg_5__3_ ( .D(n21415), .CK(clk), .QN(n18902) );
  DFF_X1 bvector3_reg_5__4_ ( .D(n21414), .CK(clk), .QN(n18939) );
  DFF_X1 bvector3_reg_5__5_ ( .D(n21413), .CK(clk), .QN(n18976) );
  DFF_X1 bvector3_reg_5__6_ ( .D(n21412), .CK(clk), .QN(n19013) );
  DFF_X1 bvector3_reg_5__7_ ( .D(n21411), .CK(clk), .QN(n19050) );
  DFF_X1 bvector3_reg_5__8_ ( .D(n21410), .CK(clk), .QN(n19087) );
  DFF_X1 bvector3_reg_5__9_ ( .D(n21409), .CK(clk), .QN(n19124) );
  DFF_X1 bvector3_reg_5__10_ ( .D(n21408), .CK(clk), .QN(n19161) );
  DFF_X1 bvector3_reg_5__11_ ( .D(n21407), .CK(clk), .QN(n19198) );
  DFF_X1 bvector3_reg_5__12_ ( .D(n21406), .CK(clk), .QN(n19235) );
  DFF_X1 bvector3_reg_5__13_ ( .D(n21405), .CK(clk), .QN(n19272) );
  DFF_X1 bvector3_reg_5__14_ ( .D(n21404), .CK(clk), .QN(n19309) );
  DFF_X1 bvector3_reg_5__15_ ( .D(n21403), .CK(clk), .QN(n19346) );
  DFF_X1 bvector3_reg_4__0_ ( .D(n21402), .CK(clk), .QN(n18790) );
  DFF_X1 bvector3_reg_4__1_ ( .D(n21401), .CK(clk), .QN(n18827) );
  DFF_X1 bvector3_reg_4__2_ ( .D(n21400), .CK(clk), .QN(n18864) );
  DFF_X1 bvector3_reg_4__3_ ( .D(n21399), .CK(clk), .QN(n18901) );
  DFF_X1 bvector3_reg_4__4_ ( .D(n21398), .CK(clk), .QN(n18938) );
  DFF_X1 bvector3_reg_4__5_ ( .D(n21397), .CK(clk), .QN(n18975) );
  DFF_X1 bvector3_reg_4__6_ ( .D(n21396), .CK(clk), .QN(n19012) );
  DFF_X1 bvector3_reg_4__7_ ( .D(n21395), .CK(clk), .QN(n19049) );
  DFF_X1 bvector3_reg_4__8_ ( .D(n21394), .CK(clk), .QN(n19086) );
  DFF_X1 bvector3_reg_4__9_ ( .D(n21393), .CK(clk), .QN(n19123) );
  DFF_X1 bvector3_reg_4__10_ ( .D(n21392), .CK(clk), .QN(n19160) );
  DFF_X1 bvector3_reg_4__11_ ( .D(n21391), .CK(clk), .QN(n19197) );
  DFF_X1 bvector3_reg_4__12_ ( .D(n21390), .CK(clk), .QN(n19234) );
  DFF_X1 bvector3_reg_4__13_ ( .D(n21389), .CK(clk), .QN(n19271) );
  DFF_X1 bvector3_reg_4__14_ ( .D(n21388), .CK(clk), .QN(n19308) );
  DFF_X1 bvector3_reg_4__15_ ( .D(n21387), .CK(clk), .QN(n19345) );
  DFF_X1 bvector3_reg_3__0_ ( .D(n21386), .CK(clk), .QN(n18786) );
  DFF_X1 bvector3_reg_3__1_ ( .D(n21385), .CK(clk), .QN(n18823) );
  DFF_X1 bvector3_reg_3__2_ ( .D(n21384), .CK(clk), .QN(n18860) );
  DFF_X1 bvector3_reg_3__3_ ( .D(n21383), .CK(clk), .QN(n18897) );
  DFF_X1 bvector3_reg_3__4_ ( .D(n21382), .CK(clk), .QN(n18934) );
  DFF_X1 bvector3_reg_3__5_ ( .D(n21381), .CK(clk), .QN(n18971) );
  DFF_X1 bvector3_reg_3__6_ ( .D(n21380), .CK(clk), .QN(n19008) );
  DFF_X1 bvector3_reg_3__7_ ( .D(n21379), .CK(clk), .QN(n19045) );
  DFF_X1 bvector3_reg_3__8_ ( .D(n21378), .CK(clk), .QN(n19082) );
  DFF_X1 bvector3_reg_3__9_ ( .D(n21377), .CK(clk), .QN(n19119) );
  DFF_X1 bvector3_reg_3__10_ ( .D(n21376), .CK(clk), .QN(n19156) );
  DFF_X1 bvector3_reg_3__11_ ( .D(n21375), .CK(clk), .QN(n19193) );
  DFF_X1 bvector3_reg_3__12_ ( .D(n21374), .CK(clk), .QN(n19230) );
  DFF_X1 bvector3_reg_3__13_ ( .D(n21373), .CK(clk), .QN(n19267) );
  DFF_X1 bvector3_reg_3__14_ ( .D(n21372), .CK(clk), .QN(n19304) );
  DFF_X1 bvector3_reg_3__15_ ( .D(n21371), .CK(clk), .QN(n19341) );
  DFF_X1 bvector3_reg_2__0_ ( .D(n21370), .CK(clk), .QN(n18785) );
  DFF_X1 bvector3_reg_2__1_ ( .D(n21369), .CK(clk), .QN(n18822) );
  DFF_X1 bvector3_reg_2__2_ ( .D(n21368), .CK(clk), .QN(n18859) );
  DFF_X1 bvector3_reg_2__3_ ( .D(n21367), .CK(clk), .QN(n18896) );
  DFF_X1 bvector3_reg_2__4_ ( .D(n21366), .CK(clk), .QN(n18933) );
  DFF_X1 bvector3_reg_2__5_ ( .D(n21365), .CK(clk), .QN(n18970) );
  DFF_X1 bvector3_reg_2__6_ ( .D(n21364), .CK(clk), .QN(n19007) );
  DFF_X1 bvector3_reg_2__7_ ( .D(n21363), .CK(clk), .QN(n19044) );
  DFF_X1 bvector3_reg_2__8_ ( .D(n21362), .CK(clk), .QN(n19081) );
  DFF_X1 bvector3_reg_2__9_ ( .D(n21361), .CK(clk), .QN(n19118) );
  DFF_X1 bvector3_reg_2__10_ ( .D(n21360), .CK(clk), .QN(n19155) );
  DFF_X1 bvector3_reg_2__11_ ( .D(n21359), .CK(clk), .QN(n19192) );
  DFF_X1 bvector3_reg_2__12_ ( .D(n21358), .CK(clk), .QN(n19229) );
  DFF_X1 bvector3_reg_2__13_ ( .D(n21357), .CK(clk), .QN(n19266) );
  DFF_X1 bvector3_reg_2__14_ ( .D(n21356), .CK(clk), .QN(n19303) );
  DFF_X1 bvector3_reg_2__15_ ( .D(n21355), .CK(clk), .QN(n19340) );
  DFF_X1 bvector0_reg_5__0_ ( .D(n21354), .CK(clk), .Q(n25699), .QN(n18782) );
  DFF_X1 bvector0_reg_5__1_ ( .D(n21353), .CK(clk), .Q(n25267), .QN(n18819) );
  DFF_X1 bvector0_reg_5__2_ ( .D(n21352), .CK(clk), .Q(n25701), .QN(n18856) );
  DFF_X1 bvector0_reg_5__3_ ( .D(n21351), .CK(clk), .Q(n25271), .QN(n18893) );
  DFF_X1 bvector0_reg_5__4_ ( .D(n21350), .CK(clk), .Q(n25703), .QN(n18930) );
  DFF_X1 bvector0_reg_5__5_ ( .D(n21349), .CK(clk), .Q(n25705), .QN(n18967) );
  DFF_X1 bvector0_reg_5__6_ ( .D(n21348), .CK(clk), .Q(n25707), .QN(n19004) );
  DFF_X1 bvector0_reg_5__7_ ( .D(n21347), .CK(clk), .Q(n25275), .QN(n19041) );
  DFF_X1 bvector0_reg_5__8_ ( .D(n21346), .CK(clk), .Q(n25709), .QN(n19078) );
  DFF_X1 bvector0_reg_5__9_ ( .D(n21345), .CK(clk), .Q(n25711), .QN(n19115) );
  DFF_X1 bvector0_reg_5__10_ ( .D(n21344), .CK(clk), .Q(n25713), .QN(n19152)
         );
  DFF_X1 bvector0_reg_5__11_ ( .D(n21343), .CK(clk), .Q(n25715), .QN(n19189)
         );
  DFF_X1 bvector0_reg_5__12_ ( .D(n21342), .CK(clk), .Q(n25717), .QN(n19226)
         );
  DFF_X1 bvector0_reg_5__13_ ( .D(n21341), .CK(clk), .Q(n25721), .QN(n19263)
         );
  DFF_X1 bvector0_reg_5__14_ ( .D(n21340), .CK(clk), .Q(n25725), .QN(n19300)
         );
  DFF_X1 bvector0_reg_5__15_ ( .D(n21339), .CK(clk), .Q(n25729), .QN(n19337)
         );
  DFF_X1 bvector0_reg_4__0_ ( .D(n21338), .CK(clk), .Q(n25212), .QN(n18781) );
  DFF_X1 bvector0_reg_4__1_ ( .D(n21337), .CK(clk), .Q(n24900), .QN(n18818) );
  DFF_X1 bvector0_reg_4__2_ ( .D(n21336), .CK(clk), .Q(n25214), .QN(n18855) );
  DFF_X1 bvector0_reg_4__3_ ( .D(n21335), .CK(clk), .Q(n24904), .QN(n18892) );
  DFF_X1 bvector0_reg_4__4_ ( .D(n21334), .CK(clk), .Q(n25216), .QN(n18929) );
  DFF_X1 bvector0_reg_4__5_ ( .D(n21333), .CK(clk), .Q(n25218), .QN(n18966) );
  DFF_X1 bvector0_reg_4__6_ ( .D(n21332), .CK(clk), .Q(n25220), .QN(n19003) );
  DFF_X1 bvector0_reg_4__7_ ( .D(n21331), .CK(clk), .Q(n24908), .QN(n19040) );
  DFF_X1 bvector0_reg_4__8_ ( .D(n21330), .CK(clk), .Q(n25222), .QN(n19077) );
  DFF_X1 bvector0_reg_4__9_ ( .D(n21329), .CK(clk), .Q(n25224), .QN(n19114) );
  DFF_X1 bvector0_reg_4__10_ ( .D(n21328), .CK(clk), .Q(n25226), .QN(n19151)
         );
  DFF_X1 bvector0_reg_4__11_ ( .D(n21327), .CK(clk), .Q(n25228), .QN(n19188)
         );
  DFF_X1 bvector0_reg_4__12_ ( .D(n21326), .CK(clk), .Q(n25230), .QN(n19225)
         );
  DFF_X1 bvector0_reg_4__13_ ( .D(n21325), .CK(clk), .Q(n25234), .QN(n19262)
         );
  DFF_X1 bvector0_reg_4__14_ ( .D(n21324), .CK(clk), .Q(n25238), .QN(n19299)
         );
  DFF_X1 bvector0_reg_4__15_ ( .D(n21323), .CK(clk), .Q(n25242), .QN(n19336)
         );
  DFF_X1 bvector0_reg_3__0_ ( .D(n21322), .CK(clk), .Q(n25054), .QN(n18777) );
  DFF_X1 bvector0_reg_3__1_ ( .D(n21321), .CK(clk), .Q(n25269), .QN(n18814) );
  DFF_X1 bvector0_reg_3__2_ ( .D(n21320), .CK(clk), .Q(n25056), .QN(n18851) );
  DFF_X1 bvector0_reg_3__3_ ( .D(n21319), .CK(clk), .Q(n25273), .QN(n18888) );
  DFF_X1 bvector0_reg_3__4_ ( .D(n21318), .CK(clk), .Q(n25058), .QN(n18925) );
  DFF_X1 bvector0_reg_3__5_ ( .D(n21317), .CK(clk), .Q(n25060), .QN(n18962) );
  DFF_X1 bvector0_reg_3__6_ ( .D(n21316), .CK(clk), .Q(n25062), .QN(n18999) );
  DFF_X1 bvector0_reg_3__7_ ( .D(n21315), .CK(clk), .Q(n25277), .QN(n19036) );
  DFF_X1 bvector0_reg_3__8_ ( .D(n21314), .CK(clk), .Q(n25064), .QN(n19073) );
  DFF_X1 bvector0_reg_3__9_ ( .D(n21313), .CK(clk), .Q(n25066), .QN(n19110) );
  DFF_X1 bvector0_reg_3__10_ ( .D(n21312), .CK(clk), .Q(n25068), .QN(n19147)
         );
  DFF_X1 bvector0_reg_3__11_ ( .D(n21311), .CK(clk), .Q(n25070), .QN(n19184)
         );
  DFF_X1 bvector0_reg_3__12_ ( .D(n21310), .CK(clk), .Q(n25719), .QN(n19221)
         );
  DFF_X1 bvector0_reg_3__13_ ( .D(n21309), .CK(clk), .Q(n25723), .QN(n19258)
         );
  DFF_X1 bvector0_reg_3__14_ ( .D(n21308), .CK(clk), .Q(n25727), .QN(n19295)
         );
  DFF_X1 bvector0_reg_3__15_ ( .D(n21307), .CK(clk), .Q(n25731), .QN(n19332)
         );
  DFF_X1 bvector0_reg_2__0_ ( .D(n21306), .CK(clk), .Q(n25053), .QN(n18776) );
  DFF_X1 bvector0_reg_2__1_ ( .D(n21305), .CK(clk), .Q(n25268), .QN(n18813) );
  DFF_X1 bvector0_reg_2__2_ ( .D(n21304), .CK(clk), .Q(n25055), .QN(n18850) );
  DFF_X1 bvector0_reg_2__3_ ( .D(n21303), .CK(clk), .Q(n25272), .QN(n18887) );
  DFF_X1 bvector0_reg_2__4_ ( .D(n21302), .CK(clk), .Q(n25057), .QN(n18924) );
  DFF_X1 bvector0_reg_2__5_ ( .D(n21301), .CK(clk), .Q(n25059), .QN(n18961) );
  DFF_X1 bvector0_reg_2__6_ ( .D(n21300), .CK(clk), .Q(n25061), .QN(n18998) );
  DFF_X1 bvector0_reg_2__7_ ( .D(n21299), .CK(clk), .Q(n25276), .QN(n19035) );
  DFF_X1 bvector0_reg_2__8_ ( .D(n21298), .CK(clk), .Q(n25063), .QN(n19072) );
  DFF_X1 bvector0_reg_2__9_ ( .D(n21297), .CK(clk), .Q(n25065), .QN(n19109) );
  DFF_X1 bvector0_reg_2__10_ ( .D(n21296), .CK(clk), .Q(n25067), .QN(n19146)
         );
  DFF_X1 bvector0_reg_2__11_ ( .D(n21295), .CK(clk), .Q(n25069), .QN(n19183)
         );
  DFF_X1 bvector0_reg_2__12_ ( .D(n21294), .CK(clk), .Q(n25718), .QN(n19220)
         );
  DFF_X1 bvector0_reg_2__13_ ( .D(n21293), .CK(clk), .Q(n25722), .QN(n19257)
         );
  DFF_X1 bvector0_reg_2__14_ ( .D(n21292), .CK(clk), .Q(n25726), .QN(n19294)
         );
  DFF_X1 bvector0_reg_2__15_ ( .D(n21291), .CK(clk), .Q(n25730), .QN(n19331)
         );
  DFF_X2 bvector0_reg_1__4_ ( .D(n23323), .CK(clk), .QN(n27946) );
  DFF_X2 bvector0_reg_1__5_ ( .D(n23324), .CK(clk), .QN(n27947) );
  DFF_X2 bvector0_reg_1__6_ ( .D(n23325), .CK(clk), .QN(n27948) );
  DFF_X2 bvector0_reg_1__7_ ( .D(n23326), .CK(clk), .QN(n27949) );
  DFF_X2 bvector0_reg_1__8_ ( .D(n23327), .CK(clk), .QN(n27950) );
  DFF_X2 bvector0_reg_1__9_ ( .D(n23328), .CK(clk), .QN(n27951) );
  DFF_X2 bvector0_reg_1__10_ ( .D(n23329), .CK(clk), .QN(n27952) );
  DFF_X2 bvector0_reg_1__11_ ( .D(n23330), .CK(clk), .QN(n27953) );
  DFF_X2 bvector0_reg_1__12_ ( .D(n23331), .CK(clk), .QN(n27954) );
  DFF_X2 bvector0_reg_0__4_ ( .D(n23339), .CK(clk), .QN(n27962) );
  DFF_X2 bvector0_reg_0__5_ ( .D(n23340), .CK(clk), .QN(n27963) );
  DFF_X2 bvector0_reg_0__6_ ( .D(n23341), .CK(clk), .QN(n27964) );
  DFF_X2 bvector0_reg_0__7_ ( .D(n23342), .CK(clk), .QN(n27965) );
  DFF_X2 bvector0_reg_0__8_ ( .D(n23343), .CK(clk), .QN(n27966) );
  DFF_X2 bvector0_reg_0__9_ ( .D(n23344), .CK(clk), .QN(n27967) );
  DFF_X2 bvector0_reg_0__10_ ( .D(n23345), .CK(clk), .QN(n27968) );
  DFF_X2 bvector0_reg_0__11_ ( .D(n23346), .CK(clk), .QN(n27969) );
  DFF_X2 bvector0_reg_0__12_ ( .D(n23347), .CK(clk), .QN(n27970) );
  DFF_X2 bvector0_reg_0__13_ ( .D(n23348), .CK(clk), .QN(n27971) );
  DFF_X2 bvector0_reg_0__14_ ( .D(n23349), .CK(clk), .QN(n27972) );
  DFF_X2 bvector0_reg_0__15_ ( .D(n23350), .CK(clk), .QN(n27973) );
  DFF_X1 bvector1_reg_5__0_ ( .D(n21290), .CK(clk), .QN(n18773) );
  DFF_X1 bvector1_reg_5__1_ ( .D(n21289), .CK(clk), .QN(n18810) );
  DFF_X1 bvector1_reg_5__2_ ( .D(n21288), .CK(clk), .QN(n18847) );
  DFF_X1 bvector1_reg_5__3_ ( .D(n21287), .CK(clk), .QN(n18884) );
  DFF_X1 bvector1_reg_5__4_ ( .D(n21286), .CK(clk), .QN(n18921) );
  DFF_X1 bvector1_reg_5__5_ ( .D(n21285), .CK(clk), .QN(n18958) );
  DFF_X1 bvector1_reg_5__6_ ( .D(n21284), .CK(clk), .QN(n18995) );
  DFF_X1 bvector1_reg_5__7_ ( .D(n21283), .CK(clk), .QN(n19032) );
  DFF_X1 bvector1_reg_5__8_ ( .D(n21282), .CK(clk), .QN(n19069) );
  DFF_X1 bvector1_reg_5__9_ ( .D(n21281), .CK(clk), .QN(n19106) );
  DFF_X1 bvector1_reg_5__10_ ( .D(n21280), .CK(clk), .QN(n19143) );
  DFF_X1 bvector1_reg_5__11_ ( .D(n21279), .CK(clk), .QN(n19180) );
  DFF_X1 bvector1_reg_5__12_ ( .D(n21278), .CK(clk), .QN(n19217) );
  DFF_X1 bvector1_reg_5__13_ ( .D(n21277), .CK(clk), .QN(n19254) );
  DFF_X1 bvector1_reg_5__14_ ( .D(n21276), .CK(clk), .QN(n19291) );
  DFF_X1 bvector1_reg_5__15_ ( .D(n21275), .CK(clk), .QN(n19328) );
  DFF_X1 bvector1_reg_4__0_ ( .D(n21274), .CK(clk), .QN(n18772) );
  DFF_X1 bvector1_reg_4__1_ ( .D(n21273), .CK(clk), .QN(n18809) );
  DFF_X1 bvector1_reg_4__2_ ( .D(n21272), .CK(clk), .QN(n18846) );
  DFF_X1 bvector1_reg_4__3_ ( .D(n21271), .CK(clk), .QN(n18883) );
  DFF_X1 bvector1_reg_4__4_ ( .D(n21270), .CK(clk), .QN(n18920) );
  DFF_X1 bvector1_reg_4__5_ ( .D(n21269), .CK(clk), .QN(n18957) );
  DFF_X1 bvector1_reg_4__6_ ( .D(n21268), .CK(clk), .QN(n18994) );
  DFF_X1 bvector1_reg_4__7_ ( .D(n21267), .CK(clk), .QN(n19031) );
  DFF_X1 bvector1_reg_4__8_ ( .D(n21266), .CK(clk), .QN(n19068) );
  DFF_X1 bvector1_reg_4__9_ ( .D(n21265), .CK(clk), .QN(n19105) );
  DFF_X1 bvector1_reg_4__10_ ( .D(n21264), .CK(clk), .QN(n19142) );
  DFF_X1 bvector1_reg_4__11_ ( .D(n21263), .CK(clk), .QN(n19179) );
  DFF_X1 bvector1_reg_4__12_ ( .D(n21262), .CK(clk), .QN(n19216) );
  DFF_X1 bvector1_reg_4__13_ ( .D(n21261), .CK(clk), .QN(n19253) );
  DFF_X1 bvector1_reg_4__14_ ( .D(n21260), .CK(clk), .QN(n19290) );
  DFF_X1 bvector1_reg_4__15_ ( .D(n21259), .CK(clk), .QN(n19327) );
  DFF_X1 bvector1_reg_3__0_ ( .D(n21258), .CK(clk), .Q(n25553), .QN(n18768) );
  DFF_X1 bvector1_reg_3__1_ ( .D(n21257), .CK(clk), .Q(n24902), .QN(n18805) );
  DFF_X1 bvector1_reg_3__2_ ( .D(n21256), .CK(clk), .Q(n25555), .QN(n18842) );
  DFF_X1 bvector1_reg_3__3_ ( .D(n21255), .CK(clk), .Q(n24906), .QN(n18879) );
  DFF_X1 bvector1_reg_3__4_ ( .D(n21254), .CK(clk), .Q(n25557), .QN(n18916) );
  DFF_X1 bvector1_reg_3__5_ ( .D(n21253), .CK(clk), .Q(n25559), .QN(n18953) );
  DFF_X1 bvector1_reg_3__6_ ( .D(n21252), .CK(clk), .Q(n25561), .QN(n18990) );
  DFF_X1 bvector1_reg_3__7_ ( .D(n21251), .CK(clk), .Q(n24910), .QN(n19027) );
  DFF_X1 bvector1_reg_3__8_ ( .D(n21250), .CK(clk), .Q(n25563), .QN(n19064) );
  DFF_X1 bvector1_reg_3__9_ ( .D(n21249), .CK(clk), .Q(n25565), .QN(n19101) );
  DFF_X1 bvector1_reg_3__10_ ( .D(n21248), .CK(clk), .Q(n25567), .QN(n19138)
         );
  DFF_X1 bvector1_reg_3__11_ ( .D(n21247), .CK(clk), .Q(n25569), .QN(n19175)
         );
  DFF_X1 bvector1_reg_3__12_ ( .D(n21246), .CK(clk), .Q(n25232), .QN(n19212)
         );
  DFF_X1 bvector1_reg_3__13_ ( .D(n21245), .CK(clk), .Q(n25236), .QN(n19249)
         );
  DFF_X1 bvector1_reg_3__14_ ( .D(n21244), .CK(clk), .Q(n25240), .QN(n19286)
         );
  DFF_X1 bvector1_reg_3__15_ ( .D(n21243), .CK(clk), .Q(n25244), .QN(n19323)
         );
  DFF_X1 bvector1_reg_2__0_ ( .D(n21242), .CK(clk), .Q(n25552), .QN(n18767) );
  DFF_X1 bvector1_reg_2__1_ ( .D(n21241), .CK(clk), .Q(n24901), .QN(n18804) );
  DFF_X1 bvector1_reg_2__2_ ( .D(n21240), .CK(clk), .Q(n25554), .QN(n18841) );
  DFF_X1 bvector1_reg_2__3_ ( .D(n21239), .CK(clk), .Q(n24905), .QN(n18878) );
  DFF_X1 bvector1_reg_2__4_ ( .D(n21238), .CK(clk), .Q(n25556), .QN(n18915) );
  DFF_X1 bvector1_reg_2__5_ ( .D(n21237), .CK(clk), .Q(n25558), .QN(n18952) );
  DFF_X1 bvector1_reg_2__6_ ( .D(n21236), .CK(clk), .Q(n25560), .QN(n18989) );
  DFF_X1 bvector1_reg_2__7_ ( .D(n21235), .CK(clk), .Q(n24909), .QN(n19026) );
  DFF_X1 bvector1_reg_2__8_ ( .D(n21234), .CK(clk), .Q(n25562), .QN(n19063) );
  DFF_X1 bvector1_reg_2__9_ ( .D(n21233), .CK(clk), .Q(n25564), .QN(n19100) );
  DFF_X1 bvector1_reg_2__10_ ( .D(n21232), .CK(clk), .Q(n25566), .QN(n19137)
         );
  DFF_X1 bvector1_reg_2__11_ ( .D(n21231), .CK(clk), .Q(n25568), .QN(n19174)
         );
  DFF_X1 bvector1_reg_2__12_ ( .D(n21230), .CK(clk), .Q(n25231), .QN(n19211)
         );
  DFF_X1 bvector1_reg_2__13_ ( .D(n21229), .CK(clk), .Q(n25235), .QN(n19248)
         );
  DFF_X1 bvector1_reg_2__14_ ( .D(n21228), .CK(clk), .Q(n25239), .QN(n19285)
         );
  DFF_X1 bvector1_reg_2__15_ ( .D(n21227), .CK(clk), .Q(n25243), .QN(n19322)
         );
  DFF_X1 bvector2_reg_5__0_ ( .D(n21226), .CK(clk), .Q(n25698), .QN(n18764) );
  DFF_X1 bvector2_reg_5__1_ ( .D(n21225), .CK(clk), .Q(n25266), .QN(n18801) );
  DFF_X1 bvector2_reg_5__2_ ( .D(n21224), .CK(clk), .Q(n25700), .QN(n18838) );
  DFF_X1 bvector2_reg_5__3_ ( .D(n21223), .CK(clk), .Q(n25270), .QN(n18875) );
  DFF_X1 bvector2_reg_5__4_ ( .D(n21222), .CK(clk), .Q(n25702), .QN(n18912) );
  DFF_X1 bvector2_reg_5__5_ ( .D(n21221), .CK(clk), .Q(n25704), .QN(n18949) );
  DFF_X1 bvector2_reg_5__6_ ( .D(n21220), .CK(clk), .Q(n25706), .QN(n18986) );
  DFF_X1 bvector2_reg_5__7_ ( .D(n21219), .CK(clk), .Q(n25274), .QN(n19023) );
  DFF_X1 bvector2_reg_5__8_ ( .D(n21218), .CK(clk), .Q(n25708), .QN(n19060) );
  DFF_X1 bvector2_reg_5__9_ ( .D(n21217), .CK(clk), .Q(n25710), .QN(n19097) );
  DFF_X1 bvector2_reg_5__10_ ( .D(n21216), .CK(clk), .Q(n25712), .QN(n19134)
         );
  DFF_X1 bvector2_reg_5__11_ ( .D(n21215), .CK(clk), .Q(n25714), .QN(n19171)
         );
  DFF_X1 bvector2_reg_5__12_ ( .D(n21214), .CK(clk), .Q(n25716), .QN(n19208)
         );
  DFF_X1 bvector2_reg_5__13_ ( .D(n21213), .CK(clk), .Q(n25720), .QN(n19245)
         );
  DFF_X1 bvector2_reg_5__14_ ( .D(n21212), .CK(clk), .Q(n25724), .QN(n19282)
         );
  DFF_X1 bvector2_reg_5__15_ ( .D(n21211), .CK(clk), .Q(n25728), .QN(n19319)
         );
  DFF_X1 bvector2_reg_4__0_ ( .D(n21210), .CK(clk), .Q(n25211), .QN(n18763) );
  DFF_X1 bvector2_reg_4__1_ ( .D(n21209), .CK(clk), .Q(n24899), .QN(n18800) );
  DFF_X1 bvector2_reg_4__2_ ( .D(n21208), .CK(clk), .Q(n25213), .QN(n18837) );
  DFF_X1 bvector2_reg_4__3_ ( .D(n21207), .CK(clk), .Q(n24903), .QN(n18874) );
  DFF_X1 bvector2_reg_4__4_ ( .D(n21206), .CK(clk), .Q(n25215), .QN(n18911) );
  DFF_X1 bvector2_reg_4__5_ ( .D(n21205), .CK(clk), .Q(n25217), .QN(n18948) );
  DFF_X1 bvector2_reg_4__6_ ( .D(n21204), .CK(clk), .Q(n25219), .QN(n18985) );
  DFF_X1 bvector2_reg_4__7_ ( .D(n21203), .CK(clk), .Q(n24907), .QN(n19022) );
  DFF_X1 bvector2_reg_4__8_ ( .D(n21202), .CK(clk), .Q(n25221), .QN(n19059) );
  DFF_X1 bvector2_reg_4__9_ ( .D(n21201), .CK(clk), .Q(n25223), .QN(n19096) );
  DFF_X1 bvector2_reg_4__10_ ( .D(n21200), .CK(clk), .Q(n25225), .QN(n19133)
         );
  DFF_X1 bvector2_reg_4__11_ ( .D(n21199), .CK(clk), .Q(n25227), .QN(n19170)
         );
  DFF_X1 bvector2_reg_4__12_ ( .D(n21198), .CK(clk), .Q(n25229), .QN(n19207)
         );
  DFF_X1 bvector2_reg_4__13_ ( .D(n21197), .CK(clk), .Q(n25233), .QN(n19244)
         );
  DFF_X1 bvector2_reg_4__14_ ( .D(n21196), .CK(clk), .Q(n25237), .QN(n19281)
         );
  DFF_X1 bvector2_reg_4__15_ ( .D(n21195), .CK(clk), .Q(n25241), .QN(n19318)
         );
  DFF_X1 bvector2_reg_3__0_ ( .D(n21194), .CK(clk), .QN(n18759) );
  DFF_X1 bvector2_reg_3__1_ ( .D(n21193), .CK(clk), .QN(n18796) );
  DFF_X1 bvector2_reg_3__2_ ( .D(n21192), .CK(clk), .QN(n18833) );
  DFF_X1 bvector2_reg_3__3_ ( .D(n21191), .CK(clk), .QN(n18870) );
  DFF_X1 bvector2_reg_3__4_ ( .D(n21190), .CK(clk), .QN(n18907) );
  DFF_X1 bvector2_reg_3__5_ ( .D(n21189), .CK(clk), .QN(n18944) );
  DFF_X1 bvector2_reg_3__6_ ( .D(n21188), .CK(clk), .QN(n18981) );
  DFF_X1 bvector2_reg_3__7_ ( .D(n21187), .CK(clk), .QN(n19018) );
  DFF_X1 bvector2_reg_3__8_ ( .D(n21186), .CK(clk), .QN(n19055) );
  DFF_X1 bvector2_reg_3__9_ ( .D(n21185), .CK(clk), .QN(n19092) );
  DFF_X1 bvector2_reg_3__10_ ( .D(n21184), .CK(clk), .QN(n19129) );
  DFF_X1 bvector2_reg_3__11_ ( .D(n21183), .CK(clk), .QN(n19166) );
  DFF_X1 bvector2_reg_3__12_ ( .D(n21182), .CK(clk), .QN(n19203) );
  DFF_X1 bvector2_reg_3__13_ ( .D(n21181), .CK(clk), .QN(n19240) );
  DFF_X1 bvector2_reg_3__14_ ( .D(n21180), .CK(clk), .QN(n19277) );
  DFF_X1 bvector2_reg_3__15_ ( .D(n21179), .CK(clk), .QN(n19314) );
  DFF_X1 bvector2_reg_2__0_ ( .D(n21178), .CK(clk), .QN(n18758) );
  DFF_X1 bvector2_reg_2__1_ ( .D(n21177), .CK(clk), .QN(n18795) );
  DFF_X1 bvector2_reg_2__2_ ( .D(n21176), .CK(clk), .QN(n18832) );
  DFF_X1 bvector2_reg_2__3_ ( .D(n21175), .CK(clk), .QN(n18869) );
  DFF_X1 bvector2_reg_2__4_ ( .D(n21174), .CK(clk), .QN(n18906) );
  DFF_X1 bvector2_reg_2__5_ ( .D(n21173), .CK(clk), .QN(n18943) );
  DFF_X1 bvector2_reg_2__6_ ( .D(n21172), .CK(clk), .QN(n18980) );
  DFF_X1 bvector2_reg_2__7_ ( .D(n21171), .CK(clk), .QN(n19017) );
  DFF_X1 bvector2_reg_2__8_ ( .D(n21170), .CK(clk), .QN(n19054) );
  DFF_X1 bvector2_reg_2__9_ ( .D(n21169), .CK(clk), .QN(n19091) );
  DFF_X1 bvector2_reg_2__10_ ( .D(n21168), .CK(clk), .QN(n19128) );
  DFF_X1 bvector2_reg_2__11_ ( .D(n21167), .CK(clk), .QN(n19165) );
  DFF_X1 bvector2_reg_2__12_ ( .D(n21166), .CK(clk), .QN(n19202) );
  DFF_X1 bvector2_reg_2__13_ ( .D(n21165), .CK(clk), .QN(n19239) );
  DFF_X1 bvector2_reg_2__14_ ( .D(n21164), .CK(clk), .QN(n19276) );
  DFF_X1 bvector2_reg_2__15_ ( .D(n21163), .CK(clk), .QN(n19313) );
  DFF_X2 dut__bvm__address_reg_6_ ( .D(n23270), .CK(clk), .Q(
        dut__bvm__address[6]), .QN(n22425) );
  DFF_X1 mac_a0_reg_0_ ( .D(n23452), .CK(clk), .Q(n4952), .QN(n18742) );
  DFF_X1 mac_a0_reg_1_ ( .D(n23453), .CK(clk), .Q(n4953), .QN(n18705) );
  DFF_X1 mac_a0_reg_2_ ( .D(n23454), .CK(clk), .Q(n4954), .QN(n18668) );
  DFF_X1 mac_a0_reg_3_ ( .D(n23455), .CK(clk), .Q(n4955), .QN(n18631) );
  DFF_X1 mac_a0_reg_4_ ( .D(n23456), .CK(clk), .Q(n4956), .QN(n18594) );
  DFF_X1 mac_a0_reg_5_ ( .D(n23457), .CK(clk), .Q(n4957), .QN(n18557) );
  DFF_X1 mac_a0_reg_6_ ( .D(n23458), .CK(clk), .Q(n4958), .QN(n18520) );
  DFF_X1 z_reg_37__0_ ( .D(n20940), .CK(clk), .Q(n25278), .QN(n20502) );
  DFF_X1 z_reg_36__0_ ( .D(n21068), .CK(clk), .QN(n20501) );
  DFF_X1 z_reg_33__0_ ( .D(n20844), .CK(clk), .QN(n20500) );
  DFF_X1 z_reg_32__0_ ( .D(n20716), .CK(clk), .QN(n20499) );
  DFF_X1 z_reg_4__0_ ( .D(n20972), .CK(clk), .QN(n20517) );
  DFF_X1 z_reg_1__0_ ( .D(n20748), .CK(clk), .QN(n20516) );
  DFF_X1 z_reg_5__0_ ( .D(n20876), .CK(clk), .Q(n25279), .QN(n20518) );
  DFF_X1 z_reg_0__0_ ( .D(n20620), .CK(clk), .QN(n20515) );
  DFF_X1 z_reg_37__1_ ( .D(n20941), .CK(clk), .Q(n25281), .QN(n20436) );
  DFF_X1 z_reg_36__1_ ( .D(n21069), .CK(clk), .QN(n20435) );
  DFF_X1 z_reg_33__1_ ( .D(n20845), .CK(clk), .QN(n20434) );
  DFF_X1 z_reg_32__1_ ( .D(n20717), .CK(clk), .QN(n20433) );
  DFF_X1 z_reg_4__1_ ( .D(n20973), .CK(clk), .QN(n20451) );
  DFF_X1 z_reg_1__1_ ( .D(n20749), .CK(clk), .QN(n20450) );
  DFF_X1 z_reg_5__1_ ( .D(n20877), .CK(clk), .Q(n25282), .QN(n20452) );
  DFF_X1 z_reg_0__1_ ( .D(n20621), .CK(clk), .QN(n20449) );
  DFF_X1 z_reg_37__2_ ( .D(n20942), .CK(clk), .Q(n25284), .QN(n20371) );
  DFF_X1 z_reg_36__2_ ( .D(n21070), .CK(clk), .QN(n20370) );
  DFF_X1 z_reg_33__2_ ( .D(n20846), .CK(clk), .QN(n20369) );
  DFF_X1 z_reg_32__2_ ( .D(n20718), .CK(clk), .QN(n20368) );
  DFF_X1 z_reg_4__2_ ( .D(n20974), .CK(clk), .QN(n20386) );
  DFF_X1 z_reg_1__2_ ( .D(n20750), .CK(clk), .QN(n20385) );
  DFF_X1 z_reg_5__2_ ( .D(n20878), .CK(clk), .Q(n25285), .QN(n20387) );
  DFF_X1 z_reg_0__2_ ( .D(n20622), .CK(clk), .QN(n20384) );
  DFF_X1 z_reg_37__3_ ( .D(n20943), .CK(clk), .Q(n25287), .QN(n20306) );
  DFF_X1 z_reg_36__3_ ( .D(n21071), .CK(clk), .QN(n20305) );
  DFF_X1 z_reg_33__3_ ( .D(n20847), .CK(clk), .QN(n20304) );
  DFF_X1 z_reg_32__3_ ( .D(n20719), .CK(clk), .QN(n20303) );
  DFF_X1 z_reg_4__3_ ( .D(n20975), .CK(clk), .QN(n20321) );
  DFF_X1 z_reg_1__3_ ( .D(n20751), .CK(clk), .QN(n20320) );
  DFF_X1 z_reg_5__3_ ( .D(n20879), .CK(clk), .Q(n25288), .QN(n20322) );
  DFF_X1 z_reg_0__3_ ( .D(n20623), .CK(clk), .QN(n20319) );
  DFF_X1 z_reg_37__4_ ( .D(n20944), .CK(clk), .Q(n25291), .QN(n20241) );
  DFF_X1 z_reg_36__4_ ( .D(n21072), .CK(clk), .QN(n20240) );
  DFF_X1 z_reg_33__4_ ( .D(n20848), .CK(clk), .QN(n20239) );
  DFF_X1 z_reg_32__4_ ( .D(n20720), .CK(clk), .QN(n20238) );
  DFF_X1 z_reg_4__4_ ( .D(n20976), .CK(clk), .QN(n20256) );
  DFF_X1 z_reg_1__4_ ( .D(n20752), .CK(clk), .QN(n20255) );
  DFF_X1 z_reg_5__4_ ( .D(n20880), .CK(clk), .Q(n25293), .QN(n20257) );
  DFF_X1 z_reg_0__4_ ( .D(n20624), .CK(clk), .QN(n20254) );
  DFF_X1 z_reg_37__5_ ( .D(n20945), .CK(clk), .Q(n25297), .QN(n20176) );
  DFF_X1 z_reg_36__5_ ( .D(n21073), .CK(clk), .QN(n20175) );
  DFF_X1 z_reg_33__5_ ( .D(n20849), .CK(clk), .QN(n20174) );
  DFF_X1 z_reg_32__5_ ( .D(n20721), .CK(clk), .QN(n20173) );
  DFF_X1 z_reg_4__5_ ( .D(n20977), .CK(clk), .QN(n20191) );
  DFF_X1 z_reg_1__5_ ( .D(n20753), .CK(clk), .QN(n20190) );
  DFF_X1 z_reg_5__5_ ( .D(n20881), .CK(clk), .Q(n25299), .QN(n20192) );
  DFF_X1 z_reg_0__5_ ( .D(n20625), .CK(clk), .QN(n20189) );
  DFF_X1 z_reg_37__6_ ( .D(n20946), .CK(clk), .Q(n25302), .QN(n20111) );
  DFF_X1 z_reg_36__6_ ( .D(n21074), .CK(clk), .QN(n20110) );
  DFF_X1 z_reg_33__6_ ( .D(n20850), .CK(clk), .QN(n20109) );
  DFF_X1 z_reg_32__6_ ( .D(n20722), .CK(clk), .QN(n20108) );
  DFF_X1 z_reg_4__6_ ( .D(n20978), .CK(clk), .QN(n20126) );
  DFF_X1 z_reg_1__6_ ( .D(n20754), .CK(clk), .QN(n20125) );
  DFF_X1 z_reg_5__6_ ( .D(n20882), .CK(clk), .Q(n25304), .QN(n20127) );
  DFF_X1 z_reg_0__6_ ( .D(n20626), .CK(clk), .QN(n20124) );
  DFF_X1 z_reg_37__7_ ( .D(n20947), .CK(clk), .Q(n25307), .QN(n20046) );
  DFF_X1 z_reg_36__7_ ( .D(n21075), .CK(clk), .QN(n20045) );
  DFF_X1 z_reg_33__7_ ( .D(n20851), .CK(clk), .QN(n20044) );
  DFF_X1 z_reg_32__7_ ( .D(n20723), .CK(clk), .QN(n20043) );
  DFF_X1 z_reg_4__7_ ( .D(n20979), .CK(clk), .QN(n20061) );
  DFF_X1 z_reg_1__7_ ( .D(n20755), .CK(clk), .QN(n20060) );
  DFF_X1 z_reg_5__7_ ( .D(n20883), .CK(clk), .Q(n25309), .QN(n20062) );
  DFF_X1 z_reg_0__7_ ( .D(n20627), .CK(clk), .QN(n20059) );
  DFF_X1 z_reg_37__8_ ( .D(n20948), .CK(clk), .Q(n25312), .QN(n19981) );
  DFF_X1 z_reg_36__8_ ( .D(n21076), .CK(clk), .QN(n19980) );
  DFF_X1 z_reg_33__8_ ( .D(n20852), .CK(clk), .QN(n19979) );
  DFF_X1 z_reg_32__8_ ( .D(n20724), .CK(clk), .QN(n19978) );
  DFF_X1 z_reg_4__8_ ( .D(n20980), .CK(clk), .QN(n19996) );
  DFF_X1 z_reg_1__8_ ( .D(n20756), .CK(clk), .QN(n19995) );
  DFF_X1 z_reg_5__8_ ( .D(n20884), .CK(clk), .Q(n25314), .QN(n19997) );
  DFF_X1 z_reg_0__8_ ( .D(n20628), .CK(clk), .QN(n19994) );
  DFF_X1 z_reg_37__9_ ( .D(n20949), .CK(clk), .Q(n25317), .QN(n19916) );
  DFF_X1 z_reg_36__9_ ( .D(n21077), .CK(clk), .QN(n19915) );
  DFF_X1 z_reg_33__9_ ( .D(n20853), .CK(clk), .QN(n19914) );
  DFF_X1 z_reg_32__9_ ( .D(n20725), .CK(clk), .QN(n19913) );
  DFF_X1 z_reg_4__9_ ( .D(n20981), .CK(clk), .QN(n19931) );
  DFF_X1 z_reg_1__9_ ( .D(n20757), .CK(clk), .QN(n19930) );
  DFF_X1 z_reg_5__9_ ( .D(n20885), .CK(clk), .Q(n25319), .QN(n19932) );
  DFF_X1 z_reg_0__9_ ( .D(n20629), .CK(clk), .QN(n19929) );
  DFF_X1 z_reg_37__10_ ( .D(n20950), .CK(clk), .Q(n25322), .QN(n19851) );
  DFF_X1 z_reg_36__10_ ( .D(n21078), .CK(clk), .QN(n19850) );
  DFF_X1 z_reg_33__10_ ( .D(n20854), .CK(clk), .QN(n19849) );
  DFF_X1 z_reg_32__10_ ( .D(n20726), .CK(clk), .QN(n19848) );
  DFF_X1 z_reg_4__10_ ( .D(n20982), .CK(clk), .QN(n19866) );
  DFF_X1 z_reg_1__10_ ( .D(n20758), .CK(clk), .QN(n19865) );
  DFF_X1 z_reg_5__10_ ( .D(n20886), .CK(clk), .Q(n25324), .QN(n19867) );
  DFF_X1 z_reg_0__10_ ( .D(n20630), .CK(clk), .QN(n19864) );
  DFF_X1 z_reg_37__11_ ( .D(n20951), .CK(clk), .Q(n25327), .QN(n19786) );
  DFF_X1 z_reg_36__11_ ( .D(n21079), .CK(clk), .QN(n19785) );
  DFF_X1 z_reg_33__11_ ( .D(n20855), .CK(clk), .QN(n19784) );
  DFF_X1 z_reg_32__11_ ( .D(n20727), .CK(clk), .QN(n19783) );
  DFF_X1 z_reg_4__11_ ( .D(n20983), .CK(clk), .QN(n19801) );
  DFF_X1 z_reg_1__11_ ( .D(n20759), .CK(clk), .QN(n19800) );
  DFF_X1 z_reg_5__11_ ( .D(n20887), .CK(clk), .Q(n25329), .QN(n19802) );
  DFF_X1 z_reg_0__11_ ( .D(n20631), .CK(clk), .QN(n19799) );
  DFF_X1 z_reg_37__12_ ( .D(n20952), .CK(clk), .Q(n25332), .QN(n19721) );
  DFF_X1 z_reg_36__12_ ( .D(n21080), .CK(clk), .QN(n19720) );
  DFF_X1 z_reg_33__12_ ( .D(n20856), .CK(clk), .QN(n19719) );
  DFF_X1 z_reg_32__12_ ( .D(n20728), .CK(clk), .QN(n19718) );
  DFF_X1 z_reg_4__12_ ( .D(n20984), .CK(clk), .QN(n19736) );
  DFF_X1 z_reg_1__12_ ( .D(n20760), .CK(clk), .QN(n19735) );
  DFF_X1 z_reg_5__12_ ( .D(n20888), .CK(clk), .Q(n25334), .QN(n19737) );
  DFF_X1 z_reg_0__12_ ( .D(n20632), .CK(clk), .QN(n19734) );
  DFF_X1 z_reg_37__13_ ( .D(n20953), .CK(clk), .Q(n25337), .QN(n19656) );
  DFF_X1 z_reg_36__13_ ( .D(n21081), .CK(clk), .QN(n19655) );
  DFF_X1 z_reg_33__13_ ( .D(n20857), .CK(clk), .QN(n19654) );
  DFF_X1 z_reg_32__13_ ( .D(n20729), .CK(clk), .QN(n19653) );
  DFF_X1 z_reg_4__13_ ( .D(n20985), .CK(clk), .QN(n19671) );
  DFF_X1 z_reg_1__13_ ( .D(n20761), .CK(clk), .QN(n19670) );
  DFF_X1 z_reg_5__13_ ( .D(n20889), .CK(clk), .Q(n25339), .QN(n19672) );
  DFF_X1 z_reg_0__13_ ( .D(n20633), .CK(clk), .QN(n19669) );
  DFF_X1 z_reg_37__14_ ( .D(n20954), .CK(clk), .Q(n25342), .QN(n19591) );
  DFF_X1 z_reg_36__14_ ( .D(n21082), .CK(clk), .QN(n19590) );
  DFF_X1 z_reg_33__14_ ( .D(n20858), .CK(clk), .QN(n19589) );
  DFF_X1 z_reg_32__14_ ( .D(n20730), .CK(clk), .QN(n19588) );
  DFF_X1 z_reg_4__14_ ( .D(n20986), .CK(clk), .QN(n19606) );
  DFF_X1 z_reg_1__14_ ( .D(n20762), .CK(clk), .QN(n19605) );
  DFF_X1 z_reg_5__14_ ( .D(n20890), .CK(clk), .Q(n25344), .QN(n19607) );
  DFF_X1 z_reg_0__14_ ( .D(n20634), .CK(clk), .QN(n19604) );
  DFF_X1 mac_a1_reg_10_ ( .D(n23478), .CK(clk), .Q(n4946), .QN(n17780) );
  DFF_X1 mac_a1_reg_11_ ( .D(n23479), .CK(clk), .Q(n4947), .QN(n17743) );
  DFF_X1 z_reg_23__0_ ( .D(n20908), .CK(clk), .Q(n25280), .QN(n20510) );
  DFF_X1 z_reg_22__0_ ( .D(n21036), .CK(clk), .QN(n20509) );
  DFF_X1 z_reg_19__0_ ( .D(n20812), .CK(clk), .QN(n20508) );
  DFF_X1 z_reg_18__0_ ( .D(n20684), .CK(clk), .QN(n20507) );
  DFF_X1 z_reg_54__0_ ( .D(n21004), .CK(clk), .QN(n20493) );
  DFF_X1 z_reg_51__0_ ( .D(n20780), .CK(clk), .QN(n20492) );
  DFF_X1 z_reg_50__0_ ( .D(n20652), .CK(clk), .Q(n25570), .QN(n20491) );
  DFF_X1 z_reg_55__0_ ( .D(n20588), .CK(clk), .Q(n25347), .QN(n20494) );
  DFF_X1 z_reg_23__1_ ( .D(n20909), .CK(clk), .Q(n25283), .QN(n20444) );
  DFF_X1 z_reg_22__1_ ( .D(n21037), .CK(clk), .QN(n20443) );
  DFF_X1 z_reg_19__1_ ( .D(n20813), .CK(clk), .QN(n20442) );
  DFF_X1 z_reg_18__1_ ( .D(n20685), .CK(clk), .QN(n20441) );
  DFF_X1 z_reg_54__1_ ( .D(n21005), .CK(clk), .QN(n20427) );
  DFF_X1 z_reg_51__1_ ( .D(n20781), .CK(clk), .QN(n20426) );
  DFF_X1 z_reg_50__1_ ( .D(n20653), .CK(clk), .Q(n25263), .QN(n20425) );
  DFF_X1 z_reg_55__1_ ( .D(n20589), .CK(clk), .Q(n25348), .QN(n20428) );
  DFF_X1 z_reg_23__2_ ( .D(n20910), .CK(clk), .Q(n25286), .QN(n20379) );
  DFF_X1 z_reg_22__2_ ( .D(n21038), .CK(clk), .QN(n20378) );
  DFF_X1 z_reg_19__2_ ( .D(n20814), .CK(clk), .QN(n20377) );
  DFF_X1 z_reg_18__2_ ( .D(n20686), .CK(clk), .QN(n20376) );
  DFF_X1 z_reg_54__2_ ( .D(n21006), .CK(clk), .QN(n20362) );
  DFF_X1 z_reg_51__2_ ( .D(n20782), .CK(clk), .QN(n20361) );
  DFF_X1 z_reg_50__2_ ( .D(n20654), .CK(clk), .Q(n25571), .QN(n20360) );
  DFF_X1 z_reg_55__2_ ( .D(n20590), .CK(clk), .Q(n25349), .QN(n20363) );
  DFF_X1 z_reg_23__3_ ( .D(n20911), .CK(clk), .Q(n25289), .QN(n20314) );
  DFF_X1 z_reg_22__3_ ( .D(n21039), .CK(clk), .QN(n20313) );
  DFF_X1 z_reg_19__3_ ( .D(n20815), .CK(clk), .QN(n20312) );
  DFF_X1 z_reg_18__3_ ( .D(n20687), .CK(clk), .QN(n20311) );
  DFF_X1 z_reg_54__3_ ( .D(n21007), .CK(clk), .QN(n20297) );
  DFF_X1 z_reg_51__3_ ( .D(n20783), .CK(clk), .QN(n20296) );
  DFF_X1 z_reg_50__3_ ( .D(n20655), .CK(clk), .Q(n25572), .QN(n20295) );
  DFF_X1 z_reg_55__3_ ( .D(n20591), .CK(clk), .Q(n25350), .QN(n20298) );
  DFF_X1 z_reg_23__4_ ( .D(n20912), .CK(clk), .Q(n25295), .QN(n20249) );
  DFF_X1 z_reg_22__4_ ( .D(n21040), .CK(clk), .QN(n20248) );
  DFF_X1 z_reg_19__4_ ( .D(n20816), .CK(clk), .QN(n20247) );
  DFF_X1 z_reg_18__4_ ( .D(n20688), .CK(clk), .QN(n20246) );
  DFF_X1 z_reg_54__4_ ( .D(n21008), .CK(clk), .QN(n20232) );
  DFF_X1 z_reg_51__4_ ( .D(n20784), .CK(clk), .QN(n20231) );
  DFF_X1 z_reg_50__4_ ( .D(n20656), .CK(clk), .Q(n25573), .QN(n20230) );
  DFF_X1 z_reg_55__4_ ( .D(n20592), .CK(clk), .Q(n25351), .QN(n20233) );
  DFF_X1 z_reg_23__5_ ( .D(n20913), .CK(clk), .Q(n25301), .QN(n20184) );
  DFF_X1 z_reg_22__5_ ( .D(n21041), .CK(clk), .QN(n20183) );
  DFF_X1 z_reg_19__5_ ( .D(n20817), .CK(clk), .QN(n20182) );
  DFF_X1 z_reg_18__5_ ( .D(n20689), .CK(clk), .QN(n20181) );
  DFF_X1 z_reg_54__5_ ( .D(n21009), .CK(clk), .QN(n20167) );
  DFF_X1 z_reg_51__5_ ( .D(n20785), .CK(clk), .QN(n20166) );
  DFF_X1 z_reg_50__5_ ( .D(n20657), .CK(clk), .Q(n25264), .QN(n20165) );
  DFF_X1 z_reg_55__5_ ( .D(n20593), .CK(clk), .Q(n25352), .QN(n20168) );
  DFF_X1 z_reg_23__6_ ( .D(n20914), .CK(clk), .Q(n25306), .QN(n20119) );
  DFF_X1 z_reg_22__6_ ( .D(n21042), .CK(clk), .QN(n20118) );
  DFF_X1 z_reg_19__6_ ( .D(n20818), .CK(clk), .QN(n20117) );
  DFF_X1 z_reg_18__6_ ( .D(n20690), .CK(clk), .QN(n20116) );
  DFF_X1 z_reg_54__6_ ( .D(n21010), .CK(clk), .QN(n20102) );
  DFF_X1 z_reg_51__6_ ( .D(n20786), .CK(clk), .QN(n20101) );
  DFF_X1 z_reg_50__6_ ( .D(n20658), .CK(clk), .Q(n25574), .QN(n20100) );
  DFF_X1 z_reg_55__6_ ( .D(n20594), .CK(clk), .Q(n25353), .QN(n20103) );
  DFF_X1 z_reg_23__7_ ( .D(n20915), .CK(clk), .Q(n25311), .QN(n20054) );
  DFF_X1 z_reg_22__7_ ( .D(n21043), .CK(clk), .QN(n20053) );
  DFF_X1 z_reg_19__7_ ( .D(n20819), .CK(clk), .QN(n20052) );
  DFF_X1 z_reg_18__7_ ( .D(n20691), .CK(clk), .QN(n20051) );
  DFF_X1 z_reg_51__7_ ( .D(n20787), .CK(clk), .QN(n20036) );
  DFF_X1 z_reg_50__7_ ( .D(n20659), .CK(clk), .Q(n25576), .QN(n20035) );
  DFF_X1 z_reg_55__7_ ( .D(n20595), .CK(clk), .Q(n25354), .QN(n20038) );
  DFF_X1 z_reg_23__8_ ( .D(n20916), .CK(clk), .Q(n25316), .QN(n19989) );
  DFF_X1 z_reg_22__8_ ( .D(n21044), .CK(clk), .QN(n19988) );
  DFF_X1 z_reg_19__8_ ( .D(n20820), .CK(clk), .QN(n19987) );
  DFF_X1 z_reg_18__8_ ( .D(n20692), .CK(clk), .QN(n19986) );
  DFF_X1 z_reg_51__8_ ( .D(n20788), .CK(clk), .QN(n19971) );
  DFF_X1 z_reg_50__8_ ( .D(n20660), .CK(clk), .Q(n25578), .QN(n19970) );
  DFF_X1 z_reg_55__8_ ( .D(n20596), .CK(clk), .Q(n25355), .QN(n19973) );
  DFF_X1 z_reg_23__9_ ( .D(n20917), .CK(clk), .Q(n25321), .QN(n19924) );
  DFF_X1 z_reg_22__9_ ( .D(n21045), .CK(clk), .QN(n19923) );
  DFF_X1 z_reg_19__9_ ( .D(n20821), .CK(clk), .QN(n19922) );
  DFF_X1 z_reg_18__9_ ( .D(n20693), .CK(clk), .QN(n19921) );
  DFF_X1 z_reg_51__9_ ( .D(n20789), .CK(clk), .QN(n19906) );
  DFF_X1 z_reg_50__9_ ( .D(n20661), .CK(clk), .Q(n25580), .QN(n19905) );
  DFF_X1 z_reg_55__9_ ( .D(n20597), .CK(clk), .Q(n25356), .QN(n19908) );
  DFF_X1 z_reg_23__10_ ( .D(n20918), .CK(clk), .Q(n25326), .QN(n19859) );
  DFF_X1 z_reg_22__10_ ( .D(n21046), .CK(clk), .QN(n19858) );
  DFF_X1 z_reg_19__10_ ( .D(n20822), .CK(clk), .QN(n19857) );
  DFF_X1 z_reg_18__10_ ( .D(n20694), .CK(clk), .QN(n19856) );
  DFF_X1 z_reg_51__10_ ( .D(n20790), .CK(clk), .QN(n19841) );
  DFF_X1 z_reg_50__10_ ( .D(n20662), .CK(clk), .Q(n25582), .QN(n19840) );
  DFF_X1 z_reg_55__10_ ( .D(n20598), .CK(clk), .Q(n25357), .QN(n19843) );
  DFF_X1 z_reg_23__11_ ( .D(n20919), .CK(clk), .Q(n25331), .QN(n19794) );
  DFF_X1 z_reg_22__11_ ( .D(n21047), .CK(clk), .QN(n19793) );
  DFF_X1 z_reg_19__11_ ( .D(n20823), .CK(clk), .QN(n19792) );
  DFF_X1 z_reg_18__11_ ( .D(n20695), .CK(clk), .QN(n19791) );
  DFF_X1 z_reg_51__11_ ( .D(n20791), .CK(clk), .QN(n19776) );
  DFF_X1 z_reg_50__11_ ( .D(n20663), .CK(clk), .Q(n25584), .QN(n19775) );
  DFF_X1 z_reg_55__11_ ( .D(n20599), .CK(clk), .Q(n25358), .QN(n19778) );
  DFF_X1 z_reg_23__12_ ( .D(n20920), .CK(clk), .Q(n25336), .QN(n19729) );
  DFF_X1 z_reg_22__12_ ( .D(n21048), .CK(clk), .QN(n19728) );
  DFF_X1 z_reg_19__12_ ( .D(n20824), .CK(clk), .QN(n19727) );
  DFF_X1 z_reg_18__12_ ( .D(n20696), .CK(clk), .QN(n19726) );
  DFF_X1 z_reg_51__12_ ( .D(n20792), .CK(clk), .QN(n19711) );
  DFF_X1 z_reg_50__12_ ( .D(n20664), .CK(clk), .Q(n25586), .QN(n19710) );
  DFF_X1 z_reg_55__12_ ( .D(n20600), .CK(clk), .Q(n25359), .QN(n19713) );
  DFF_X1 z_reg_23__13_ ( .D(n20921), .CK(clk), .Q(n25341), .QN(n19664) );
  DFF_X1 z_reg_22__13_ ( .D(n21049), .CK(clk), .QN(n19663) );
  DFF_X1 z_reg_19__13_ ( .D(n20825), .CK(clk), .QN(n19662) );
  DFF_X1 z_reg_18__13_ ( .D(n20697), .CK(clk), .QN(n19661) );
  DFF_X1 z_reg_51__13_ ( .D(n20793), .CK(clk), .QN(n19646) );
  DFF_X1 z_reg_50__13_ ( .D(n20665), .CK(clk), .Q(n25588), .QN(n19645) );
  DFF_X1 z_reg_55__13_ ( .D(n20601), .CK(clk), .Q(n25360), .QN(n19648) );
  DFF_X1 z_reg_23__14_ ( .D(n20922), .CK(clk), .Q(n25346), .QN(n19599) );
  DFF_X1 z_reg_22__14_ ( .D(n21050), .CK(clk), .QN(n19598) );
  DFF_X1 z_reg_19__14_ ( .D(n20826), .CK(clk), .QN(n19597) );
  DFF_X1 z_reg_18__14_ ( .D(n20698), .CK(clk), .QN(n19596) );
  DFF_X1 z_reg_51__14_ ( .D(n20794), .CK(clk), .QN(n19581) );
  DFF_X1 z_reg_50__14_ ( .D(n20666), .CK(clk), .Q(n25590), .QN(n19580) );
  DFF_X1 mac_a2_reg_0_ ( .D(n23484), .CK(clk), .Q(n4920), .QN(n17558) );
  DFF_X1 mac_a2_reg_1_ ( .D(n23485), .CK(clk), .Q(n4921), .QN(n17521) );
  DFF_X1 mac_a2_reg_2_ ( .D(n23486), .CK(clk), .Q(n4922), .QN(n17484) );
  DFF_X1 mac_a2_reg_3_ ( .D(n23487), .CK(clk), .Q(n4923), .QN(n17447) );
  DFF_X1 mac_a2_reg_4_ ( .D(n23488), .CK(clk), .Q(n4924), .QN(n17410) );
  DFF_X1 mac_a2_reg_5_ ( .D(n23489), .CK(clk), .Q(n4925), .QN(n17373) );
  DFF_X1 mac_a2_reg_6_ ( .D(n23490), .CK(clk), .Q(n4926), .QN(n17336) );
  DFF_X1 mac_a2_reg_7_ ( .D(n23491), .CK(clk), .Q(n4927), .QN(n17299) );
  DFF_X1 mac_a2_reg_8_ ( .D(n23492), .CK(clk), .Q(n4928), .QN(n17262) );
  DFF_X1 mac_a2_reg_9_ ( .D(n23493), .CK(clk), .Q(n4929), .QN(n17225) );
  DFF_X1 mac_a2_reg_10_ ( .D(n23494), .CK(clk), .Q(n4930), .QN(n17188) );
  DFF_X1 mac_a2_reg_11_ ( .D(n23495), .CK(clk), .Q(n4931), .QN(n17151) );
  DFF_X1 z_reg_61__1_ ( .D(n20573), .CK(clk), .QN(n20432) );
  DFF_X1 z_reg_61__2_ ( .D(n20574), .CK(clk), .QN(n20367) );
  DFF_X1 z_reg_61__3_ ( .D(n20575), .CK(clk), .QN(n20302) );
  DFF_X1 z_reg_45__4_ ( .D(n20928), .CK(clk), .QN(n20245) );
  DFF_X1 z_reg_44__4_ ( .D(n21056), .CK(clk), .Q(n24911), .QN(n20244) );
  DFF_X1 z_reg_41__4_ ( .D(n20832), .CK(clk), .Q(n25290), .QN(n20243) );
  DFF_X1 z_reg_40__4_ ( .D(n20704), .CK(clk), .Q(n24912), .QN(n20242) );
  DFF_X1 z_reg_12__4_ ( .D(n20960), .CK(clk), .QN(n20260) );
  DFF_X1 z_reg_9__4_ ( .D(n20736), .CK(clk), .QN(n20259) );
  DFF_X1 z_reg_13__4_ ( .D(n20864), .CK(clk), .Q(n25292), .QN(n20261) );
  DFF_X1 z_reg_8__4_ ( .D(n20608), .CK(clk), .Q(n24914), .QN(n20258) );
  DFF_X1 z_reg_61__4_ ( .D(n20576), .CK(clk), .QN(n20237) );
  DFF_X1 z_reg_45__5_ ( .D(n20929), .CK(clk), .QN(n20180) );
  DFF_X1 z_reg_44__5_ ( .D(n21057), .CK(clk), .Q(n24917), .QN(n20179) );
  DFF_X1 z_reg_41__5_ ( .D(n20833), .CK(clk), .Q(n25296), .QN(n20178) );
  DFF_X1 z_reg_40__5_ ( .D(n20705), .CK(clk), .Q(n24918), .QN(n20177) );
  DFF_X1 z_reg_12__5_ ( .D(n20961), .CK(clk), .QN(n20195) );
  DFF_X1 z_reg_9__5_ ( .D(n20737), .CK(clk), .QN(n20194) );
  DFF_X1 z_reg_13__5_ ( .D(n20865), .CK(clk), .Q(n25298), .QN(n20196) );
  DFF_X1 z_reg_8__5_ ( .D(n20609), .CK(clk), .Q(n24920), .QN(n20193) );
  DFF_X1 z_reg_61__5_ ( .D(n20577), .CK(clk), .QN(n20172) );
  DFF_X1 z_reg_45__6_ ( .D(n20930), .CK(clk), .QN(n20115) );
  DFF_X1 z_reg_44__6_ ( .D(n21058), .CK(clk), .Q(n25575), .QN(n20114) );
  DFF_X1 z_reg_41__6_ ( .D(n20834), .CK(clk), .Q(n25071), .QN(n20113) );
  DFF_X1 z_reg_40__6_ ( .D(n20706), .CK(clk), .Q(n24923), .QN(n20112) );
  DFF_X1 z_reg_12__6_ ( .D(n20962), .CK(clk), .QN(n20130) );
  DFF_X1 z_reg_9__6_ ( .D(n20738), .CK(clk), .QN(n20129) );
  DFF_X1 z_reg_13__6_ ( .D(n20866), .CK(clk), .Q(n25303), .QN(n20131) );
  DFF_X1 z_reg_8__6_ ( .D(n20610), .CK(clk), .Q(n24925), .QN(n20128) );
  DFF_X1 z_reg_61__6_ ( .D(n20578), .CK(clk), .QN(n20107) );
  DFF_X1 z_reg_45__7_ ( .D(n20931), .CK(clk), .QN(n20050) );
  DFF_X1 z_reg_44__7_ ( .D(n21059), .CK(clk), .Q(n25577), .QN(n20049) );
  DFF_X1 z_reg_41__7_ ( .D(n20835), .CK(clk), .Q(n25072), .QN(n20048) );
  DFF_X1 z_reg_40__7_ ( .D(n20707), .CK(clk), .Q(n24928), .QN(n20047) );
  DFF_X1 z_reg_12__7_ ( .D(n20963), .CK(clk), .QN(n20065) );
  DFF_X1 z_reg_9__7_ ( .D(n20739), .CK(clk), .QN(n20064) );
  DFF_X1 z_reg_13__7_ ( .D(n20867), .CK(clk), .Q(n25308), .QN(n20066) );
  DFF_X1 z_reg_8__7_ ( .D(n20611), .CK(clk), .Q(n24930), .QN(n20063) );
  DFF_X1 z_reg_61__7_ ( .D(n20579), .CK(clk), .QN(n20042) );
  DFF_X1 z_reg_45__8_ ( .D(n20932), .CK(clk), .QN(n19985) );
  DFF_X1 z_reg_44__8_ ( .D(n21060), .CK(clk), .Q(n25579), .QN(n19984) );
  DFF_X1 z_reg_41__8_ ( .D(n20836), .CK(clk), .Q(n25073), .QN(n19983) );
  DFF_X1 z_reg_40__8_ ( .D(n20708), .CK(clk), .Q(n24933), .QN(n19982) );
  DFF_X1 z_reg_12__8_ ( .D(n20964), .CK(clk), .QN(n20000) );
  DFF_X1 z_reg_9__8_ ( .D(n20740), .CK(clk), .QN(n19999) );
  DFF_X1 z_reg_13__8_ ( .D(n20868), .CK(clk), .Q(n25313), .QN(n20001) );
  DFF_X1 z_reg_8__8_ ( .D(n20612), .CK(clk), .Q(n24935), .QN(n19998) );
  DFF_X1 z_reg_61__8_ ( .D(n20580), .CK(clk), .QN(n19977) );
  DFF_X1 z_reg_45__9_ ( .D(n20933), .CK(clk), .QN(n19920) );
  DFF_X1 z_reg_44__9_ ( .D(n21061), .CK(clk), .Q(n25581), .QN(n19919) );
  DFF_X1 z_reg_41__9_ ( .D(n20837), .CK(clk), .Q(n25074), .QN(n19918) );
  DFF_X1 z_reg_40__9_ ( .D(n20709), .CK(clk), .Q(n24938), .QN(n19917) );
  DFF_X1 z_reg_12__9_ ( .D(n20965), .CK(clk), .QN(n19935) );
  DFF_X1 z_reg_9__9_ ( .D(n20741), .CK(clk), .QN(n19934) );
  DFF_X1 z_reg_13__9_ ( .D(n20869), .CK(clk), .Q(n25318), .QN(n19936) );
  DFF_X1 z_reg_8__9_ ( .D(n20613), .CK(clk), .Q(n24940), .QN(n19933) );
  DFF_X1 z_reg_61__9_ ( .D(n20581), .CK(clk), .QN(n19912) );
  DFF_X1 z_reg_45__10_ ( .D(n20934), .CK(clk), .QN(n19855) );
  DFF_X1 z_reg_44__10_ ( .D(n21062), .CK(clk), .Q(n25583), .QN(n19854) );
  DFF_X1 z_reg_41__10_ ( .D(n20838), .CK(clk), .Q(n25075), .QN(n19853) );
  DFF_X1 z_reg_40__10_ ( .D(n20710), .CK(clk), .Q(n24943), .QN(n19852) );
  DFF_X1 z_reg_12__10_ ( .D(n20966), .CK(clk), .QN(n19870) );
  DFF_X1 z_reg_9__10_ ( .D(n20742), .CK(clk), .QN(n19869) );
  DFF_X1 z_reg_13__10_ ( .D(n20870), .CK(clk), .Q(n25323), .QN(n19871) );
  DFF_X1 z_reg_8__10_ ( .D(n20614), .CK(clk), .Q(n24945), .QN(n19868) );
  DFF_X1 z_reg_61__10_ ( .D(n20582), .CK(clk), .QN(n19847) );
  DFF_X1 z_reg_45__11_ ( .D(n20935), .CK(clk), .QN(n19790) );
  DFF_X1 z_reg_44__11_ ( .D(n21063), .CK(clk), .Q(n25585), .QN(n19789) );
  DFF_X1 z_reg_41__11_ ( .D(n20839), .CK(clk), .Q(n25076), .QN(n19788) );
  DFF_X1 z_reg_40__11_ ( .D(n20711), .CK(clk), .Q(n24948), .QN(n19787) );
  DFF_X1 z_reg_12__11_ ( .D(n20967), .CK(clk), .QN(n19805) );
  DFF_X1 z_reg_9__11_ ( .D(n20743), .CK(clk), .QN(n19804) );
  DFF_X1 z_reg_13__11_ ( .D(n20871), .CK(clk), .Q(n25328), .QN(n19806) );
  DFF_X1 z_reg_8__11_ ( .D(n20615), .CK(clk), .Q(n24950), .QN(n19803) );
  DFF_X1 z_reg_61__11_ ( .D(n20583), .CK(clk), .QN(n19782) );
  DFF_X1 z_reg_45__12_ ( .D(n20936), .CK(clk), .QN(n19725) );
  DFF_X1 z_reg_44__12_ ( .D(n21064), .CK(clk), .Q(n25587), .QN(n19724) );
  DFF_X1 z_reg_41__12_ ( .D(n20840), .CK(clk), .Q(n25077), .QN(n19723) );
  DFF_X1 z_reg_40__12_ ( .D(n20712), .CK(clk), .Q(n24953), .QN(n19722) );
  DFF_X1 z_reg_12__12_ ( .D(n20968), .CK(clk), .QN(n19740) );
  DFF_X1 z_reg_9__12_ ( .D(n20744), .CK(clk), .QN(n19739) );
  DFF_X1 z_reg_13__12_ ( .D(n20872), .CK(clk), .Q(n25333), .QN(n19741) );
  DFF_X1 z_reg_8__12_ ( .D(n20616), .CK(clk), .Q(n24955), .QN(n19738) );
  DFF_X1 z_reg_61__12_ ( .D(n20584), .CK(clk), .QN(n19717) );
  DFF_X1 z_reg_45__13_ ( .D(n20937), .CK(clk), .QN(n19660) );
  DFF_X1 z_reg_44__13_ ( .D(n21065), .CK(clk), .Q(n25589), .QN(n19659) );
  DFF_X1 z_reg_41__13_ ( .D(n20841), .CK(clk), .Q(n25078), .QN(n19658) );
  DFF_X1 z_reg_40__13_ ( .D(n20713), .CK(clk), .Q(n24958), .QN(n19657) );
  DFF_X1 z_reg_12__13_ ( .D(n20969), .CK(clk), .QN(n19675) );
  DFF_X1 z_reg_9__13_ ( .D(n20745), .CK(clk), .QN(n19674) );
  DFF_X1 z_reg_13__13_ ( .D(n20873), .CK(clk), .Q(n25338), .QN(n19676) );
  DFF_X1 z_reg_8__13_ ( .D(n20617), .CK(clk), .Q(n24960), .QN(n19673) );
  DFF_X1 z_reg_61__13_ ( .D(n20585), .CK(clk), .QN(n19652) );
  DFF_X1 z_reg_45__14_ ( .D(n20938), .CK(clk), .QN(n19595) );
  DFF_X1 z_reg_44__14_ ( .D(n21066), .CK(clk), .Q(n25591), .QN(n19594) );
  DFF_X1 z_reg_41__14_ ( .D(n20842), .CK(clk), .Q(n25079), .QN(n19593) );
  DFF_X1 z_reg_40__14_ ( .D(n20714), .CK(clk), .Q(n24963), .QN(n19592) );
  DFF_X1 z_reg_12__14_ ( .D(n20970), .CK(clk), .QN(n19610) );
  DFF_X1 z_reg_9__14_ ( .D(n20746), .CK(clk), .QN(n19609) );
  DFF_X1 z_reg_13__14_ ( .D(n20874), .CK(clk), .Q(n25343), .QN(n19611) );
  DFF_X1 z_reg_8__14_ ( .D(n20618), .CK(clk), .Q(n24964), .QN(n19608) );
  DFF_X1 z_reg_61__14_ ( .D(n20586), .CK(clk), .QN(n19587) );
  DFF_X1 mac_a3_reg_6_ ( .D(n23506), .CK(clk), .Q(n4910), .QN(n16744) );
  DFF_X1 mac_a3_reg_8_ ( .D(n23508), .CK(clk), .Q(n4912), .QN(n16670) );
  DFF_X1 mac_a3_reg_9_ ( .D(n23509), .CK(clk), .Q(n4913), .QN(n16633) );
  DFF_X1 mac_a3_reg_10_ ( .D(n23510), .CK(clk), .Q(n4914), .QN(n16596) );
  DFF_X1 z_reg_31__4_ ( .D(n20896), .CK(clk), .QN(n20253) );
  DFF_X1 z_reg_30__4_ ( .D(n21024), .CK(clk), .Q(n24915), .QN(n20252) );
  DFF_X1 z_reg_27__4_ ( .D(n20800), .CK(clk), .Q(n25294), .QN(n20251) );
  DFF_X1 z_reg_26__4_ ( .D(n20672), .CK(clk), .Q(n24916), .QN(n20250) );
  DFF_X1 z_reg_58__4_ ( .D(n20640), .CK(clk), .Q(n24913), .QN(n20234) );
  DFF_X1 z_reg_31__5_ ( .D(n20897), .CK(clk), .QN(n20188) );
  DFF_X1 z_reg_30__5_ ( .D(n21025), .CK(clk), .Q(n24921), .QN(n20187) );
  DFF_X1 z_reg_27__5_ ( .D(n20801), .CK(clk), .Q(n25300), .QN(n20186) );
  DFF_X1 z_reg_26__5_ ( .D(n20673), .CK(clk), .Q(n24922), .QN(n20185) );
  DFF_X1 z_reg_58__5_ ( .D(n20641), .CK(clk), .Q(n24919), .QN(n20169) );
  DFF_X1 z_reg_31__6_ ( .D(n20898), .CK(clk), .QN(n20123) );
  DFF_X1 z_reg_30__6_ ( .D(n21026), .CK(clk), .Q(n24926), .QN(n20122) );
  DFF_X1 z_reg_27__6_ ( .D(n20802), .CK(clk), .Q(n25305), .QN(n20121) );
  DFF_X1 z_reg_26__6_ ( .D(n20674), .CK(clk), .Q(n24927), .QN(n20120) );
  DFF_X1 z_reg_58__6_ ( .D(n20642), .CK(clk), .Q(n24924), .QN(n20104) );
  DFF_X1 mac_z_reg_6_ ( .D(n20549), .CK(clk), .Q(n642), .QN(n20132) );
  DFF_X1 z_reg_31__7_ ( .D(n20899), .CK(clk), .QN(n20058) );
  DFF_X1 z_reg_30__7_ ( .D(n21027), .CK(clk), .Q(n24931), .QN(n20057) );
  DFF_X1 z_reg_27__7_ ( .D(n20803), .CK(clk), .Q(n25310), .QN(n20056) );
  DFF_X1 z_reg_26__7_ ( .D(n20675), .CK(clk), .Q(n24932), .QN(n20055) );
  DFF_X1 z_reg_58__7_ ( .D(n20643), .CK(clk), .Q(n24929), .QN(n20039) );
  DFF_X1 z_reg_31__8_ ( .D(n20900), .CK(clk), .QN(n19993) );
  DFF_X1 z_reg_30__8_ ( .D(n21028), .CK(clk), .Q(n24936), .QN(n19992) );
  DFF_X1 z_reg_27__8_ ( .D(n20804), .CK(clk), .Q(n25315), .QN(n19991) );
  DFF_X1 z_reg_26__8_ ( .D(n20676), .CK(clk), .Q(n24937), .QN(n19990) );
  DFF_X1 z_reg_58__8_ ( .D(n20644), .CK(clk), .Q(n24934), .QN(n19974) );
  DFF_X1 mac_z_reg_8_ ( .D(n20547), .CK(clk), .Q(n644), .QN(n20002) );
  DFF_X1 z_reg_31__9_ ( .D(n20901), .CK(clk), .QN(n19928) );
  DFF_X1 z_reg_30__9_ ( .D(n21029), .CK(clk), .Q(n24941), .QN(n19927) );
  DFF_X1 z_reg_27__9_ ( .D(n20805), .CK(clk), .Q(n25320), .QN(n19926) );
  DFF_X1 z_reg_26__9_ ( .D(n20677), .CK(clk), .Q(n24942), .QN(n19925) );
  DFF_X1 z_reg_58__9_ ( .D(n20645), .CK(clk), .Q(n24939), .QN(n19909) );
  DFF_X1 mac_z_reg_9_ ( .D(n20546), .CK(clk), .Q(n645), .QN(n19937) );
  DFF_X1 z_reg_31__10_ ( .D(n20902), .CK(clk), .QN(n19863) );
  DFF_X1 z_reg_30__10_ ( .D(n21030), .CK(clk), .Q(n24946), .QN(n19862) );
  DFF_X1 z_reg_27__10_ ( .D(n20806), .CK(clk), .Q(n25325), .QN(n19861) );
  DFF_X1 z_reg_26__10_ ( .D(n20678), .CK(clk), .Q(n24947), .QN(n19860) );
  DFF_X1 z_reg_58__10_ ( .D(n20646), .CK(clk), .Q(n24944), .QN(n19844) );
  DFF_X1 z_reg_31__11_ ( .D(n20903), .CK(clk), .QN(n19798) );
  DFF_X1 z_reg_30__11_ ( .D(n21031), .CK(clk), .Q(n24951), .QN(n19797) );
  DFF_X1 z_reg_27__11_ ( .D(n20807), .CK(clk), .Q(n25330), .QN(n19796) );
  DFF_X1 z_reg_26__11_ ( .D(n20679), .CK(clk), .Q(n24952), .QN(n19795) );
  DFF_X1 z_reg_58__11_ ( .D(n20647), .CK(clk), .Q(n24949), .QN(n19779) );
  DFF_X1 z_reg_31__12_ ( .D(n20904), .CK(clk), .QN(n19733) );
  DFF_X1 z_reg_30__12_ ( .D(n21032), .CK(clk), .Q(n24956), .QN(n19732) );
  DFF_X1 z_reg_27__12_ ( .D(n20808), .CK(clk), .Q(n25335), .QN(n19731) );
  DFF_X1 z_reg_26__12_ ( .D(n20680), .CK(clk), .Q(n24957), .QN(n19730) );
  DFF_X1 z_reg_58__12_ ( .D(n20648), .CK(clk), .Q(n24954), .QN(n19714) );
  DFF_X1 z_reg_31__13_ ( .D(n20905), .CK(clk), .QN(n19668) );
  DFF_X1 z_reg_30__13_ ( .D(n21033), .CK(clk), .Q(n24961), .QN(n19667) );
  DFF_X1 z_reg_27__13_ ( .D(n20809), .CK(clk), .Q(n25340), .QN(n19666) );
  DFF_X1 z_reg_26__13_ ( .D(n20681), .CK(clk), .Q(n24962), .QN(n19665) );
  DFF_X1 z_reg_58__13_ ( .D(n20649), .CK(clk), .Q(n24959), .QN(n19649) );
  DFF_X1 z_reg_31__14_ ( .D(n20906), .CK(clk), .QN(n19603) );
  DFF_X1 z_reg_30__14_ ( .D(n21034), .CK(clk), .Q(n24965), .QN(n19602) );
  DFF_X1 z_reg_27__14_ ( .D(n20810), .CK(clk), .Q(n25345), .QN(n19601) );
  DFF_X1 z_reg_26__14_ ( .D(n20682), .CK(clk), .Q(n24966), .QN(n19600) );
  DFF_X1 z_reg_58__14_ ( .D(n20650), .CK(clk), .Q(n25265), .QN(n19584) );
  AND2_X1 U833 ( .A1(n11202), .A2(n11203), .ZN(n11192) );
  AND2_X1 U849 ( .A1(n11212), .A2(n24892), .ZN(n11207) );
  AND2_X1 U879 ( .A1(n11202), .A2(n11235), .ZN(n11194) );
  AND2_X1 U882 ( .A1(n11236), .A2(n25251), .ZN(n11226) );
  AND2_X1 U885 ( .A1(n11236), .A2(n11212), .ZN(n11231) );
  AND2_X1 U898 ( .A1(n11236), .A2(n11235), .ZN(n11245) );
  AND2_X1 U900 ( .A1(n11236), .A2(n11203), .ZN(n11244) );
  AND2_X1 U912 ( .A1(n11257), .A2(n11212), .ZN(n11225) );
  AND2_X1 U915 ( .A1(n11257), .A2(n11235), .ZN(n11221) );
  AND2_X1 U917 ( .A1(n11257), .A2(n25251), .ZN(n11227) );
  AND2_X1 U930 ( .A1(n11235), .A2(n24892), .ZN(n11266) );
  AND2_X1 U933 ( .A1(n24892), .A2(n11203), .ZN(n11265) );
  AND2_X1 U948 ( .A1(n25251), .A2(n11202), .ZN(n11276) );
  AND2_X1 U952 ( .A1(n11202), .A2(n11212), .ZN(n11275) );
  AND2_X1 U1563 ( .A1(n11436), .A2(n19349), .ZN(n11433) );
  OR3_X1 U5764 ( .A1(n26295), .A2(n22406), .A3(n26283), .ZN(n13084) );
  AND2_X1 U7560 ( .A1(n22396), .A2(n22395), .ZN(n15515) );
  OR2_X1 U7599 ( .A1(n15530), .A2(n15537), .ZN(n15531) );
  AND2_X1 U10525 ( .A1(n11257), .A2(n11203), .ZN(n11220) );
  OAI22_X2 U3 ( .A1(n19547), .A2(n26130), .B1(n10080), .B2(n10081), .ZN(n20540) );
  NOR4_X2 U4 ( .A1(n10082), .A2(n10083), .A3(n10084), .A4(n10085), .ZN(n10080)
         );
  NAND4_X2 U5 ( .A1(n10086), .A2(n10087), .A3(n10088), .A4(n10089), .ZN(n10085) );
  AOI221_X2 U6 ( .B1(n10090), .B2(n26186), .C1(n10092), .C2(n26160), .A(n10094), .ZN(n10089) );
  OAI22_X2 U7 ( .A1(n19533), .A2(n10095), .B1(n19532), .B2(n10096), .ZN(n10094) );
  AOI221_X2 U10 ( .B1(n10097), .B2(n26158), .C1(n10099), .C2(n26156), .A(
        n10101), .ZN(n10088) );
  OAI22_X2 U11 ( .A1(n19539), .A2(n10102), .B1(n19538), .B2(n10103), .ZN(
        n10101) );
  AOI221_X2 U15 ( .B1(n10104), .B2(n26147), .C1(n10106), .C2(n26178), .A(
        n10108), .ZN(n10087) );
  OAI22_X2 U16 ( .A1(n19541), .A2(n10109), .B1(n19540), .B2(n10110), .ZN(
        n10108) );
  AOI221_X2 U19 ( .B1(n10111), .B2(n26174), .C1(n19490), .C2(n26139), .A(
        n10114), .ZN(n10086) );
  OAI22_X2 U20 ( .A1(n19545), .A2(n10115), .B1(n19544), .B2(n10116), .ZN(
        n10114) );
  NAND4_X2 U22 ( .A1(n10117), .A2(n10118), .A3(n10119), .A4(n10120), .ZN(
        n10084) );
  AOI221_X2 U23 ( .B1(n10121), .B2(n26191), .C1(n10123), .C2(n26161), .A(
        n10125), .ZN(n10120) );
  OAI22_X2 U24 ( .A1(n19517), .A2(n10126), .B1(n19516), .B2(n10127), .ZN(
        n10125) );
  AOI221_X2 U27 ( .B1(n10128), .B2(n26159), .C1(n10130), .C2(n26171), .A(
        n10132), .ZN(n10119) );
  OAI22_X2 U28 ( .A1(n19523), .A2(n10133), .B1(n19522), .B2(n10134), .ZN(
        n10132) );
  AOI221_X2 U31 ( .B1(n10135), .B2(n26146), .C1(n10137), .C2(n26177), .A(
        n10139), .ZN(n10118) );
  OAI22_X2 U32 ( .A1(n19525), .A2(n10140), .B1(n19524), .B2(n10141), .ZN(
        n10139) );
  AOI221_X2 U35 ( .B1(n10142), .B2(n26175), .C1(n10144), .C2(n26170), .A(
        n10146), .ZN(n10117) );
  OAI22_X2 U36 ( .A1(n19531), .A2(n10147), .B1(n19530), .B2(n10148), .ZN(
        n10146) );
  NAND4_X2 U39 ( .A1(n10149), .A2(n10150), .A3(n10151), .A4(n10152), .ZN(
        n10083) );
  AOI221_X2 U40 ( .B1(n19496), .B2(n10153), .C1(n19495), .C2(n10154), .A(
        n10155), .ZN(n10152) );
  OAI22_X2 U41 ( .A1(n10156), .A2(n28693), .B1(n10158), .B2(n28692), .ZN(
        n10155) );
  AOI221_X2 U42 ( .B1(n19492), .B2(n10160), .C1(n19491), .C2(n10161), .A(
        n10162), .ZN(n10151) );
  OAI22_X2 U43 ( .A1(n10163), .A2(n28380), .B1(n10165), .B2(n28379), .ZN(
        n10162) );
  AOI221_X2 U44 ( .B1(n19487), .B2(n10167), .C1(n19486), .C2(n10168), .A(
        n10169), .ZN(n10150) );
  OAI22_X2 U45 ( .A1(n10170), .A2(n28510), .B1(n10172), .B2(n28694), .ZN(
        n10169) );
  AOI221_X2 U46 ( .B1(n19483), .B2(n10174), .C1(n10175), .C2(n26190), .A(
        n10177), .ZN(n10149) );
  OAI22_X2 U47 ( .A1(n10178), .A2(n28257), .B1(n10180), .B2(n28256), .ZN(
        n10177) );
  NAND4_X2 U49 ( .A1(n10182), .A2(n10183), .A3(n10184), .A4(n10185), .ZN(
        n10082) );
  AOI221_X2 U50 ( .B1(n19514), .B2(n10186), .C1(n19513), .C2(n10187), .A(
        n10188), .ZN(n10185) );
  OAI22_X2 U51 ( .A1(n10189), .A2(n28696), .B1(n10191), .B2(n28695), .ZN(
        n10188) );
  AOI221_X2 U52 ( .B1(n19508), .B2(n10193), .C1(n19507), .C2(n10194), .A(
        n10195), .ZN(n10184) );
  OAI22_X2 U53 ( .A1(n10196), .A2(n28381), .B1(n10198), .B2(n28382), .ZN(
        n10195) );
  AOI221_X2 U54 ( .B1(n19504), .B2(n10200), .C1(n19503), .C2(n10201), .A(
        n10202), .ZN(n10183) );
  OAI22_X2 U55 ( .A1(n10203), .A2(n28509), .B1(n10205), .B2(n28508), .ZN(
        n10202) );
  AOI221_X2 U56 ( .B1(n19500), .B2(n10207), .C1(n19499), .C2(n10208), .A(
        n10209), .ZN(n10182) );
  OAI22_X2 U57 ( .A1(n10210), .A2(n28255), .B1(n10212), .B2(n28254), .ZN(
        n10209) );
  OAI22_X2 U58 ( .A1(n19612), .A2(n26130), .B1(n10214), .B2(n10081), .ZN(
        n20541) );
  NOR4_X2 U59 ( .A1(n10215), .A2(n10216), .A3(n10217), .A4(n10218), .ZN(n10214) );
  NAND4_X2 U60 ( .A1(n10219), .A2(n10220), .A3(n10221), .A4(n10222), .ZN(
        n10218) );
  AOI221_X2 U61 ( .B1(n10090), .B2(n25346), .C1(n10092), .C2(n24966), .A(
        n10225), .ZN(n10222) );
  OAI22_X2 U62 ( .A1(n19598), .A2(n10095), .B1(n19597), .B2(n10096), .ZN(
        n10225) );
  AOI221_X2 U65 ( .B1(n10097), .B2(n25345), .C1(n10099), .C2(n24965), .A(
        n10228), .ZN(n10221) );
  OAI22_X2 U66 ( .A1(n19604), .A2(n10102), .B1(n19603), .B2(n10103), .ZN(
        n10228) );
  AOI221_X2 U69 ( .B1(n10104), .B2(n25344), .C1(n10106), .C2(n24964), .A(
        n10231), .ZN(n10220) );
  OAI22_X2 U70 ( .A1(n19606), .A2(n10109), .B1(n19605), .B2(n10110), .ZN(
        n10231) );
  AOI221_X2 U73 ( .B1(n10111), .B2(n25343), .C1(n19555), .C2(n26139), .A(
        n10233), .ZN(n10219) );
  OAI22_X2 U74 ( .A1(n19610), .A2(n10115), .B1(n19609), .B2(n10116), .ZN(
        n10233) );
  NAND4_X2 U76 ( .A1(n10234), .A2(n10235), .A3(n10236), .A4(n10237), .ZN(
        n10217) );
  AOI221_X2 U77 ( .B1(n10121), .B2(n28378), .C1(n10123), .C2(n25265), .A(
        n10240), .ZN(n10237) );
  OAI22_X2 U78 ( .A1(n19582), .A2(n10126), .B1(n19581), .B2(n10127), .ZN(
        n10240) );
  AOI221_X2 U81 ( .B1(n10128), .B2(n28691), .C1(n10130), .C2(n28507), .A(
        n10243), .ZN(n10236) );
  OAI22_X2 U82 ( .A1(n19588), .A2(n10133), .B1(n19587), .B2(n10134), .ZN(
        n10243) );
  AOI221_X2 U85 ( .B1(n10135), .B2(n25342), .C1(n10137), .C2(n24963), .A(
        n10246), .ZN(n10235) );
  OAI22_X2 U86 ( .A1(n19590), .A2(n10140), .B1(n19589), .B2(n10141), .ZN(
        n10246) );
  AOI221_X2 U89 ( .B1(n10142), .B2(n25079), .C1(n10144), .C2(n25591), .A(
        n10249), .ZN(n10234) );
  OAI22_X2 U90 ( .A1(n19596), .A2(n10147), .B1(n19595), .B2(n10148), .ZN(
        n10249) );
  NAND4_X2 U93 ( .A1(n10250), .A2(n10251), .A3(n10252), .A4(n10253), .ZN(
        n10216) );
  AOI221_X2 U94 ( .B1(n19561), .B2(n10153), .C1(n19560), .C2(n10154), .A(
        n10254), .ZN(n10253) );
  OAI22_X2 U95 ( .A1(n10156), .A2(n28682), .B1(n10158), .B2(n28681), .ZN(
        n10254) );
  AOI221_X2 U96 ( .B1(n19557), .B2(n10160), .C1(n19556), .C2(n10161), .A(
        n10257), .ZN(n10252) );
  OAI22_X2 U97 ( .A1(n10163), .A2(n28371), .B1(n10165), .B2(n28370), .ZN(
        n10257) );
  AOI221_X2 U98 ( .B1(n19552), .B2(n10167), .C1(n19551), .C2(n10168), .A(
        n10260), .ZN(n10251) );
  OAI22_X2 U99 ( .A1(n10170), .A2(n28505), .B1(n10172), .B2(n28685), .ZN(
        n10260) );
  AOI221_X2 U100 ( .B1(n19548), .B2(n10174), .C1(n10175), .C2(n25590), .A(
        n10264), .ZN(n10250) );
  OAI22_X2 U101 ( .A1(n10178), .A2(n28251), .B1(n10180), .B2(n28250), .ZN(
        n10264) );
  NAND4_X2 U103 ( .A1(n10267), .A2(n10268), .A3(n10269), .A4(n10270), .ZN(
        n10215) );
  AOI221_X2 U104 ( .B1(n19579), .B2(n10186), .C1(n19578), .C2(n10187), .A(
        n10271), .ZN(n10270) );
  OAI22_X2 U105 ( .A1(n10189), .A2(n28689), .B1(n10191), .B2(n28687), .ZN(
        n10271) );
  AOI221_X2 U106 ( .B1(n19573), .B2(n10193), .C1(n19572), .C2(n10194), .A(
        n10274), .ZN(n10269) );
  OAI22_X2 U107 ( .A1(n10196), .A2(n28374), .B1(n10198), .B2(n28376), .ZN(
        n10274) );
  AOI221_X2 U108 ( .B1(n19569), .B2(n10200), .C1(n19568), .C2(n10201), .A(
        n10277), .ZN(n10268) );
  OAI22_X2 U109 ( .A1(n10203), .A2(n28502), .B1(n10205), .B2(n28501), .ZN(
        n10277) );
  AOI221_X2 U110 ( .B1(n19565), .B2(n10207), .C1(n19564), .C2(n10208), .A(
        n10280), .ZN(n10267) );
  OAI22_X2 U111 ( .A1(n10210), .A2(n28247), .B1(n10212), .B2(n28246), .ZN(
        n10280) );
  OAI22_X2 U112 ( .A1(n19677), .A2(n26130), .B1(n10283), .B2(n10081), .ZN(
        n20542) );
  NOR4_X2 U113 ( .A1(n10284), .A2(n10285), .A3(n10286), .A4(n10287), .ZN(
        n10283) );
  NAND4_X2 U114 ( .A1(n10288), .A2(n10289), .A3(n10290), .A4(n10291), .ZN(
        n10287) );
  AOI221_X2 U115 ( .B1(n10090), .B2(n25341), .C1(n10092), .C2(n24962), .A(
        n10294), .ZN(n10291) );
  OAI22_X2 U116 ( .A1(n19663), .A2(n10095), .B1(n19662), .B2(n10096), .ZN(
        n10294) );
  AOI221_X2 U119 ( .B1(n10097), .B2(n25340), .C1(n10099), .C2(n24961), .A(
        n10297), .ZN(n10290) );
  OAI22_X2 U120 ( .A1(n19669), .A2(n10102), .B1(n19668), .B2(n10103), .ZN(
        n10297) );
  AOI221_X2 U123 ( .B1(n10104), .B2(n25339), .C1(n10106), .C2(n24960), .A(
        n10300), .ZN(n10289) );
  OAI22_X2 U124 ( .A1(n19671), .A2(n10109), .B1(n19670), .B2(n10110), .ZN(
        n10300) );
  AOI221_X2 U127 ( .B1(n10111), .B2(n25338), .C1(n19620), .C2(n26139), .A(
        n10302), .ZN(n10288) );
  OAI22_X2 U128 ( .A1(n19675), .A2(n10115), .B1(n19674), .B2(n10116), .ZN(
        n10302) );
  NAND4_X2 U130 ( .A1(n10303), .A2(n10304), .A3(n10305), .A4(n10306), .ZN(
        n10286) );
  AOI221_X2 U131 ( .B1(n10121), .B2(n25360), .C1(n10123), .C2(n24959), .A(
        n10309), .ZN(n10306) );
  OAI22_X2 U132 ( .A1(n19647), .A2(n10126), .B1(n19646), .B2(n10127), .ZN(
        n10309) );
  AOI221_X2 U135 ( .B1(n10128), .B2(n28680), .C1(n10130), .C2(n28500), .A(
        n10312), .ZN(n10305) );
  OAI22_X2 U136 ( .A1(n19653), .A2(n10133), .B1(n19652), .B2(n10134), .ZN(
        n10312) );
  AOI221_X2 U139 ( .B1(n10135), .B2(n25337), .C1(n10137), .C2(n24958), .A(
        n10315), .ZN(n10304) );
  OAI22_X2 U140 ( .A1(n19655), .A2(n10140), .B1(n19654), .B2(n10141), .ZN(
        n10315) );
  AOI221_X2 U143 ( .B1(n10142), .B2(n25078), .C1(n10144), .C2(n25589), .A(
        n10318), .ZN(n10303) );
  OAI22_X2 U144 ( .A1(n19661), .A2(n10147), .B1(n19660), .B2(n10148), .ZN(
        n10318) );
  NAND4_X2 U147 ( .A1(n10319), .A2(n10320), .A3(n10321), .A4(n10322), .ZN(
        n10285) );
  AOI221_X2 U148 ( .B1(n19626), .B2(n10153), .C1(n19625), .C2(n10154), .A(
        n10323), .ZN(n10322) );
  OAI22_X2 U149 ( .A1(n10156), .A2(n28671), .B1(n10158), .B2(n28670), .ZN(
        n10323) );
  AOI221_X2 U150 ( .B1(n19622), .B2(n10160), .C1(n19621), .C2(n10161), .A(
        n10326), .ZN(n10321) );
  OAI22_X2 U151 ( .A1(n10163), .A2(n28363), .B1(n10165), .B2(n28362), .ZN(
        n10326) );
  AOI221_X2 U152 ( .B1(n19617), .B2(n10167), .C1(n19616), .C2(n10168), .A(
        n10329), .ZN(n10320) );
  OAI22_X2 U153 ( .A1(n10170), .A2(n28498), .B1(n10172), .B2(n28674), .ZN(
        n10329) );
  AOI221_X2 U154 ( .B1(n19613), .B2(n10174), .C1(n10175), .C2(n25588), .A(
        n10333), .ZN(n10319) );
  OAI22_X2 U155 ( .A1(n10178), .A2(n28243), .B1(n10180), .B2(n28242), .ZN(
        n10333) );
  NAND4_X2 U157 ( .A1(n10336), .A2(n10337), .A3(n10338), .A4(n10339), .ZN(
        n10284) );
  AOI221_X2 U158 ( .B1(n19644), .B2(n10186), .C1(n19643), .C2(n10187), .A(
        n10340), .ZN(n10339) );
  OAI22_X2 U159 ( .A1(n10189), .A2(n28678), .B1(n10191), .B2(n28676), .ZN(
        n10340) );
  AOI221_X2 U160 ( .B1(n19638), .B2(n10193), .C1(n19637), .C2(n10194), .A(
        n10343), .ZN(n10338) );
  OAI22_X2 U161 ( .A1(n10196), .A2(n28366), .B1(n10198), .B2(n28368), .ZN(
        n10343) );
  AOI221_X2 U162 ( .B1(n19634), .B2(n10200), .C1(n19633), .C2(n10201), .A(
        n10346), .ZN(n10337) );
  OAI22_X2 U163 ( .A1(n10203), .A2(n28495), .B1(n10205), .B2(n28494), .ZN(
        n10346) );
  AOI221_X2 U164 ( .B1(n19630), .B2(n10207), .C1(n19629), .C2(n10208), .A(
        n10349), .ZN(n10336) );
  OAI22_X2 U165 ( .A1(n10210), .A2(n28239), .B1(n10212), .B2(n28238), .ZN(
        n10349) );
  OAI22_X2 U166 ( .A1(n19742), .A2(n26130), .B1(n10352), .B2(n10081), .ZN(
        n20543) );
  NOR4_X2 U167 ( .A1(n10353), .A2(n10354), .A3(n10355), .A4(n10356), .ZN(
        n10352) );
  NAND4_X2 U168 ( .A1(n10357), .A2(n10358), .A3(n10359), .A4(n10360), .ZN(
        n10356) );
  AOI221_X2 U169 ( .B1(n10090), .B2(n25336), .C1(n10092), .C2(n24957), .A(
        n10363), .ZN(n10360) );
  OAI22_X2 U170 ( .A1(n19728), .A2(n10095), .B1(n19727), .B2(n10096), .ZN(
        n10363) );
  AOI221_X2 U173 ( .B1(n10097), .B2(n25335), .C1(n10099), .C2(n24956), .A(
        n10366), .ZN(n10359) );
  OAI22_X2 U174 ( .A1(n19734), .A2(n10102), .B1(n19733), .B2(n10103), .ZN(
        n10366) );
  AOI221_X2 U177 ( .B1(n10104), .B2(n25334), .C1(n10106), .C2(n24955), .A(
        n10369), .ZN(n10358) );
  OAI22_X2 U178 ( .A1(n19736), .A2(n10109), .B1(n19735), .B2(n10110), .ZN(
        n10369) );
  AOI221_X2 U181 ( .B1(n10111), .B2(n25333), .C1(n19685), .C2(n26139), .A(
        n10371), .ZN(n10357) );
  OAI22_X2 U182 ( .A1(n19740), .A2(n10115), .B1(n19739), .B2(n10116), .ZN(
        n10371) );
  NAND4_X2 U184 ( .A1(n10372), .A2(n10373), .A3(n10374), .A4(n10375), .ZN(
        n10355) );
  AOI221_X2 U185 ( .B1(n10121), .B2(n25359), .C1(n10123), .C2(n24954), .A(
        n10378), .ZN(n10375) );
  OAI22_X2 U186 ( .A1(n19712), .A2(n10126), .B1(n19711), .B2(n10127), .ZN(
        n10378) );
  AOI221_X2 U189 ( .B1(n10128), .B2(n28669), .C1(n10130), .C2(n28493), .A(
        n10381), .ZN(n10374) );
  OAI22_X2 U190 ( .A1(n19718), .A2(n10133), .B1(n19717), .B2(n10134), .ZN(
        n10381) );
  AOI221_X2 U193 ( .B1(n10135), .B2(n25332), .C1(n10137), .C2(n24953), .A(
        n10384), .ZN(n10373) );
  OAI22_X2 U194 ( .A1(n19720), .A2(n10140), .B1(n19719), .B2(n10141), .ZN(
        n10384) );
  AOI221_X2 U197 ( .B1(n10142), .B2(n25077), .C1(n10144), .C2(n25587), .A(
        n10387), .ZN(n10372) );
  OAI22_X2 U198 ( .A1(n19726), .A2(n10147), .B1(n19725), .B2(n10148), .ZN(
        n10387) );
  NAND4_X2 U201 ( .A1(n10388), .A2(n10389), .A3(n10390), .A4(n10391), .ZN(
        n10354) );
  AOI221_X2 U202 ( .B1(n19691), .B2(n10153), .C1(n19690), .C2(n10154), .A(
        n10392), .ZN(n10391) );
  OAI22_X2 U203 ( .A1(n10156), .A2(n28660), .B1(n10158), .B2(n28659), .ZN(
        n10392) );
  AOI221_X2 U204 ( .B1(n19687), .B2(n10160), .C1(n19686), .C2(n10161), .A(
        n10395), .ZN(n10390) );
  OAI22_X2 U205 ( .A1(n10163), .A2(n28355), .B1(n10165), .B2(n28354), .ZN(
        n10395) );
  AOI221_X2 U206 ( .B1(n19682), .B2(n10167), .C1(n19681), .C2(n10168), .A(
        n10398), .ZN(n10389) );
  OAI22_X2 U207 ( .A1(n10170), .A2(n28491), .B1(n10172), .B2(n28663), .ZN(
        n10398) );
  AOI221_X2 U208 ( .B1(n19678), .B2(n10174), .C1(n10175), .C2(n25586), .A(
        n10402), .ZN(n10388) );
  OAI22_X2 U209 ( .A1(n10178), .A2(n28235), .B1(n10180), .B2(n28234), .ZN(
        n10402) );
  NAND4_X2 U211 ( .A1(n10405), .A2(n10406), .A3(n10407), .A4(n10408), .ZN(
        n10353) );
  AOI221_X2 U212 ( .B1(n19709), .B2(n10186), .C1(n19708), .C2(n10187), .A(
        n10409), .ZN(n10408) );
  OAI22_X2 U213 ( .A1(n10189), .A2(n28667), .B1(n10191), .B2(n28665), .ZN(
        n10409) );
  AOI221_X2 U214 ( .B1(n19703), .B2(n10193), .C1(n19702), .C2(n10194), .A(
        n10412), .ZN(n10407) );
  OAI22_X2 U215 ( .A1(n10196), .A2(n28358), .B1(n10198), .B2(n28360), .ZN(
        n10412) );
  AOI221_X2 U216 ( .B1(n19699), .B2(n10200), .C1(n19698), .C2(n10201), .A(
        n10415), .ZN(n10406) );
  OAI22_X2 U217 ( .A1(n10203), .A2(n28488), .B1(n10205), .B2(n28487), .ZN(
        n10415) );
  AOI221_X2 U218 ( .B1(n19695), .B2(n10207), .C1(n19694), .C2(n10208), .A(
        n10418), .ZN(n10405) );
  OAI22_X2 U219 ( .A1(n10210), .A2(n28231), .B1(n10212), .B2(n28230), .ZN(
        n10418) );
  OAI22_X2 U220 ( .A1(n19807), .A2(n26130), .B1(n10421), .B2(n10081), .ZN(
        n20544) );
  NOR4_X2 U221 ( .A1(n10422), .A2(n10423), .A3(n10424), .A4(n10425), .ZN(
        n10421) );
  NAND4_X2 U222 ( .A1(n10426), .A2(n10427), .A3(n10428), .A4(n10429), .ZN(
        n10425) );
  AOI221_X2 U223 ( .B1(n10090), .B2(n25331), .C1(n10092), .C2(n24952), .A(
        n10432), .ZN(n10429) );
  OAI22_X2 U224 ( .A1(n19793), .A2(n10095), .B1(n19792), .B2(n10096), .ZN(
        n10432) );
  AOI221_X2 U227 ( .B1(n10097), .B2(n25330), .C1(n10099), .C2(n24951), .A(
        n10435), .ZN(n10428) );
  OAI22_X2 U228 ( .A1(n19799), .A2(n10102), .B1(n19798), .B2(n10103), .ZN(
        n10435) );
  AOI221_X2 U231 ( .B1(n10104), .B2(n25329), .C1(n10106), .C2(n24950), .A(
        n10438), .ZN(n10427) );
  OAI22_X2 U232 ( .A1(n19801), .A2(n10109), .B1(n19800), .B2(n10110), .ZN(
        n10438) );
  AOI221_X2 U235 ( .B1(n10111), .B2(n25328), .C1(n19750), .C2(n26139), .A(
        n10440), .ZN(n10426) );
  OAI22_X2 U236 ( .A1(n19805), .A2(n10115), .B1(n19804), .B2(n10116), .ZN(
        n10440) );
  NAND4_X2 U238 ( .A1(n10441), .A2(n10442), .A3(n10443), .A4(n10444), .ZN(
        n10424) );
  AOI221_X2 U239 ( .B1(n10121), .B2(n25358), .C1(n10123), .C2(n24949), .A(
        n10447), .ZN(n10444) );
  OAI22_X2 U240 ( .A1(n19777), .A2(n10126), .B1(n19776), .B2(n10127), .ZN(
        n10447) );
  AOI221_X2 U243 ( .B1(n10128), .B2(n28658), .C1(n10130), .C2(n28486), .A(
        n10450), .ZN(n10443) );
  OAI22_X2 U244 ( .A1(n19783), .A2(n10133), .B1(n19782), .B2(n10134), .ZN(
        n10450) );
  AOI221_X2 U247 ( .B1(n10135), .B2(n25327), .C1(n10137), .C2(n24948), .A(
        n10453), .ZN(n10442) );
  OAI22_X2 U248 ( .A1(n19785), .A2(n10140), .B1(n19784), .B2(n10141), .ZN(
        n10453) );
  AOI221_X2 U251 ( .B1(n10142), .B2(n25076), .C1(n10144), .C2(n25585), .A(
        n10456), .ZN(n10441) );
  OAI22_X2 U252 ( .A1(n19791), .A2(n10147), .B1(n19790), .B2(n10148), .ZN(
        n10456) );
  NAND4_X2 U255 ( .A1(n10457), .A2(n10458), .A3(n10459), .A4(n10460), .ZN(
        n10423) );
  AOI221_X2 U256 ( .B1(n19756), .B2(n10153), .C1(n19755), .C2(n10154), .A(
        n10461), .ZN(n10460) );
  OAI22_X2 U257 ( .A1(n10156), .A2(n28649), .B1(n10158), .B2(n28648), .ZN(
        n10461) );
  AOI221_X2 U258 ( .B1(n19752), .B2(n10160), .C1(n19751), .C2(n10161), .A(
        n10464), .ZN(n10459) );
  OAI22_X2 U259 ( .A1(n10163), .A2(n28347), .B1(n10165), .B2(n28346), .ZN(
        n10464) );
  AOI221_X2 U260 ( .B1(n19747), .B2(n10167), .C1(n19746), .C2(n10168), .A(
        n10467), .ZN(n10458) );
  OAI22_X2 U261 ( .A1(n10170), .A2(n28484), .B1(n10172), .B2(n28652), .ZN(
        n10467) );
  AOI221_X2 U262 ( .B1(n19743), .B2(n10174), .C1(n10175), .C2(n25584), .A(
        n10471), .ZN(n10457) );
  OAI22_X2 U263 ( .A1(n10178), .A2(n28227), .B1(n10180), .B2(n28226), .ZN(
        n10471) );
  NAND4_X2 U265 ( .A1(n10474), .A2(n10475), .A3(n10476), .A4(n10477), .ZN(
        n10422) );
  AOI221_X2 U266 ( .B1(n19774), .B2(n10186), .C1(n19773), .C2(n10187), .A(
        n10478), .ZN(n10477) );
  OAI22_X2 U267 ( .A1(n10189), .A2(n28656), .B1(n10191), .B2(n28654), .ZN(
        n10478) );
  AOI221_X2 U268 ( .B1(n19768), .B2(n10193), .C1(n19767), .C2(n10194), .A(
        n10481), .ZN(n10476) );
  OAI22_X2 U269 ( .A1(n10196), .A2(n28350), .B1(n10198), .B2(n28352), .ZN(
        n10481) );
  AOI221_X2 U270 ( .B1(n19764), .B2(n10200), .C1(n19763), .C2(n10201), .A(
        n10484), .ZN(n10475) );
  OAI22_X2 U271 ( .A1(n10203), .A2(n28481), .B1(n10205), .B2(n28480), .ZN(
        n10484) );
  AOI221_X2 U272 ( .B1(n19760), .B2(n10207), .C1(n19759), .C2(n10208), .A(
        n10487), .ZN(n10474) );
  OAI22_X2 U273 ( .A1(n10210), .A2(n28223), .B1(n10212), .B2(n28222), .ZN(
        n10487) );
  OAI22_X2 U274 ( .A1(n19872), .A2(n26130), .B1(n10490), .B2(n10081), .ZN(
        n20545) );
  NOR4_X2 U275 ( .A1(n10491), .A2(n10492), .A3(n10493), .A4(n10494), .ZN(
        n10490) );
  NAND4_X2 U276 ( .A1(n10495), .A2(n10496), .A3(n10497), .A4(n10498), .ZN(
        n10494) );
  AOI221_X2 U277 ( .B1(n10090), .B2(n25326), .C1(n10092), .C2(n24947), .A(
        n10501), .ZN(n10498) );
  OAI22_X2 U278 ( .A1(n19858), .A2(n10095), .B1(n19857), .B2(n10096), .ZN(
        n10501) );
  AOI221_X2 U281 ( .B1(n10097), .B2(n25325), .C1(n10099), .C2(n24946), .A(
        n10504), .ZN(n10497) );
  OAI22_X2 U282 ( .A1(n19864), .A2(n10102), .B1(n19863), .B2(n10103), .ZN(
        n10504) );
  AOI221_X2 U285 ( .B1(n10104), .B2(n25324), .C1(n10106), .C2(n24945), .A(
        n10507), .ZN(n10496) );
  OAI22_X2 U286 ( .A1(n19866), .A2(n10109), .B1(n19865), .B2(n10110), .ZN(
        n10507) );
  AOI221_X2 U289 ( .B1(n10111), .B2(n25323), .C1(n19815), .C2(n26139), .A(
        n10509), .ZN(n10495) );
  OAI22_X2 U290 ( .A1(n19870), .A2(n10115), .B1(n19869), .B2(n10116), .ZN(
        n10509) );
  NAND4_X2 U292 ( .A1(n10510), .A2(n10511), .A3(n10512), .A4(n10513), .ZN(
        n10493) );
  AOI221_X2 U293 ( .B1(n10121), .B2(n25357), .C1(n10123), .C2(n24944), .A(
        n10516), .ZN(n10513) );
  OAI22_X2 U294 ( .A1(n19842), .A2(n10126), .B1(n19841), .B2(n10127), .ZN(
        n10516) );
  AOI221_X2 U297 ( .B1(n10128), .B2(n28647), .C1(n10130), .C2(n28479), .A(
        n10519), .ZN(n10512) );
  OAI22_X2 U298 ( .A1(n19848), .A2(n10133), .B1(n19847), .B2(n10134), .ZN(
        n10519) );
  AOI221_X2 U301 ( .B1(n10135), .B2(n25322), .C1(n10137), .C2(n24943), .A(
        n10522), .ZN(n10511) );
  OAI22_X2 U302 ( .A1(n19850), .A2(n10140), .B1(n19849), .B2(n10141), .ZN(
        n10522) );
  AOI221_X2 U305 ( .B1(n10142), .B2(n25075), .C1(n10144), .C2(n25583), .A(
        n10525), .ZN(n10510) );
  OAI22_X2 U306 ( .A1(n19856), .A2(n10147), .B1(n19855), .B2(n10148), .ZN(
        n10525) );
  NAND4_X2 U309 ( .A1(n10526), .A2(n10527), .A3(n10528), .A4(n10529), .ZN(
        n10492) );
  AOI221_X2 U310 ( .B1(n19821), .B2(n10153), .C1(n19820), .C2(n10154), .A(
        n10530), .ZN(n10529) );
  OAI22_X2 U311 ( .A1(n10156), .A2(n28638), .B1(n10158), .B2(n28637), .ZN(
        n10530) );
  AOI221_X2 U312 ( .B1(n19817), .B2(n10160), .C1(n19816), .C2(n10161), .A(
        n10533), .ZN(n10528) );
  OAI22_X2 U313 ( .A1(n10163), .A2(n28339), .B1(n10165), .B2(n28338), .ZN(
        n10533) );
  AOI221_X2 U314 ( .B1(n19812), .B2(n10167), .C1(n19811), .C2(n10168), .A(
        n10536), .ZN(n10527) );
  OAI22_X2 U315 ( .A1(n10170), .A2(n28477), .B1(n10172), .B2(n28641), .ZN(
        n10536) );
  AOI221_X2 U316 ( .B1(n19808), .B2(n10174), .C1(n10175), .C2(n25582), .A(
        n10540), .ZN(n10526) );
  OAI22_X2 U317 ( .A1(n10178), .A2(n28219), .B1(n10180), .B2(n28218), .ZN(
        n10540) );
  NAND4_X2 U319 ( .A1(n10543), .A2(n10544), .A3(n10545), .A4(n10546), .ZN(
        n10491) );
  AOI221_X2 U320 ( .B1(n19839), .B2(n10186), .C1(n19838), .C2(n10187), .A(
        n10547), .ZN(n10546) );
  OAI22_X2 U321 ( .A1(n10189), .A2(n28645), .B1(n10191), .B2(n28643), .ZN(
        n10547) );
  AOI221_X2 U322 ( .B1(n19833), .B2(n10193), .C1(n19832), .C2(n10194), .A(
        n10550), .ZN(n10545) );
  OAI22_X2 U323 ( .A1(n10196), .A2(n28342), .B1(n10198), .B2(n28344), .ZN(
        n10550) );
  AOI221_X2 U324 ( .B1(n19829), .B2(n10200), .C1(n19828), .C2(n10201), .A(
        n10553), .ZN(n10544) );
  OAI22_X2 U325 ( .A1(n10203), .A2(n28474), .B1(n10205), .B2(n28473), .ZN(
        n10553) );
  AOI221_X2 U326 ( .B1(n19825), .B2(n10207), .C1(n19824), .C2(n10208), .A(
        n10556), .ZN(n10543) );
  OAI22_X2 U327 ( .A1(n10210), .A2(n28215), .B1(n10212), .B2(n28214), .ZN(
        n10556) );
  OAI22_X2 U328 ( .A1(n19937), .A2(n26130), .B1(n10559), .B2(n10081), .ZN(
        n20546) );
  NOR4_X2 U329 ( .A1(n10560), .A2(n10561), .A3(n10562), .A4(n10563), .ZN(
        n10559) );
  NAND4_X2 U330 ( .A1(n10564), .A2(n10565), .A3(n10566), .A4(n10567), .ZN(
        n10563) );
  AOI221_X2 U331 ( .B1(n10090), .B2(n25321), .C1(n10092), .C2(n24942), .A(
        n10570), .ZN(n10567) );
  OAI22_X2 U332 ( .A1(n19923), .A2(n10095), .B1(n19922), .B2(n10096), .ZN(
        n10570) );
  AOI221_X2 U335 ( .B1(n10097), .B2(n25320), .C1(n10099), .C2(n24941), .A(
        n10573), .ZN(n10566) );
  OAI22_X2 U336 ( .A1(n19929), .A2(n10102), .B1(n19928), .B2(n10103), .ZN(
        n10573) );
  AOI221_X2 U339 ( .B1(n10104), .B2(n25319), .C1(n10106), .C2(n24940), .A(
        n10576), .ZN(n10565) );
  OAI22_X2 U340 ( .A1(n19931), .A2(n10109), .B1(n19930), .B2(n10110), .ZN(
        n10576) );
  AOI221_X2 U343 ( .B1(n10111), .B2(n25318), .C1(n19880), .C2(n26139), .A(
        n10578), .ZN(n10564) );
  OAI22_X2 U344 ( .A1(n19935), .A2(n10115), .B1(n19934), .B2(n10116), .ZN(
        n10578) );
  NAND4_X2 U346 ( .A1(n10579), .A2(n10580), .A3(n10581), .A4(n10582), .ZN(
        n10562) );
  AOI221_X2 U347 ( .B1(n10121), .B2(n25356), .C1(n10123), .C2(n24939), .A(
        n10585), .ZN(n10582) );
  OAI22_X2 U348 ( .A1(n19907), .A2(n10126), .B1(n19906), .B2(n10127), .ZN(
        n10585) );
  AOI221_X2 U351 ( .B1(n10128), .B2(n28636), .C1(n10130), .C2(n28472), .A(
        n10588), .ZN(n10581) );
  OAI22_X2 U352 ( .A1(n19913), .A2(n10133), .B1(n19912), .B2(n10134), .ZN(
        n10588) );
  AOI221_X2 U355 ( .B1(n10135), .B2(n25317), .C1(n10137), .C2(n24938), .A(
        n10591), .ZN(n10580) );
  OAI22_X2 U356 ( .A1(n19915), .A2(n10140), .B1(n19914), .B2(n10141), .ZN(
        n10591) );
  AOI221_X2 U359 ( .B1(n10142), .B2(n25074), .C1(n10144), .C2(n25581), .A(
        n10594), .ZN(n10579) );
  OAI22_X2 U360 ( .A1(n19921), .A2(n10147), .B1(n19920), .B2(n10148), .ZN(
        n10594) );
  NAND4_X2 U363 ( .A1(n10595), .A2(n10596), .A3(n10597), .A4(n10598), .ZN(
        n10561) );
  AOI221_X2 U364 ( .B1(n19886), .B2(n10153), .C1(n19885), .C2(n10154), .A(
        n10599), .ZN(n10598) );
  OAI22_X2 U365 ( .A1(n10156), .A2(n28627), .B1(n10158), .B2(n28626), .ZN(
        n10599) );
  AOI221_X2 U366 ( .B1(n19882), .B2(n10160), .C1(n19881), .C2(n10161), .A(
        n10602), .ZN(n10597) );
  OAI22_X2 U367 ( .A1(n10163), .A2(n28331), .B1(n10165), .B2(n28330), .ZN(
        n10602) );
  AOI221_X2 U368 ( .B1(n19877), .B2(n10167), .C1(n19876), .C2(n10168), .A(
        n10605), .ZN(n10596) );
  OAI22_X2 U369 ( .A1(n10170), .A2(n28470), .B1(n10172), .B2(n28630), .ZN(
        n10605) );
  AOI221_X2 U370 ( .B1(n19873), .B2(n10174), .C1(n10175), .C2(n25580), .A(
        n10609), .ZN(n10595) );
  OAI22_X2 U371 ( .A1(n10178), .A2(n28211), .B1(n10180), .B2(n28210), .ZN(
        n10609) );
  NAND4_X2 U373 ( .A1(n10612), .A2(n10613), .A3(n10614), .A4(n10615), .ZN(
        n10560) );
  AOI221_X2 U374 ( .B1(n19904), .B2(n10186), .C1(n19903), .C2(n10187), .A(
        n10616), .ZN(n10615) );
  OAI22_X2 U375 ( .A1(n10189), .A2(n28634), .B1(n10191), .B2(n28632), .ZN(
        n10616) );
  AOI221_X2 U376 ( .B1(n19898), .B2(n10193), .C1(n19897), .C2(n10194), .A(
        n10619), .ZN(n10614) );
  OAI22_X2 U377 ( .A1(n10196), .A2(n28334), .B1(n10198), .B2(n28336), .ZN(
        n10619) );
  AOI221_X2 U378 ( .B1(n19894), .B2(n10200), .C1(n19893), .C2(n10201), .A(
        n10622), .ZN(n10613) );
  OAI22_X2 U379 ( .A1(n10203), .A2(n28467), .B1(n10205), .B2(n28466), .ZN(
        n10622) );
  AOI221_X2 U380 ( .B1(n19890), .B2(n10207), .C1(n19889), .C2(n10208), .A(
        n10625), .ZN(n10612) );
  OAI22_X2 U381 ( .A1(n10210), .A2(n28207), .B1(n10212), .B2(n28206), .ZN(
        n10625) );
  OAI22_X2 U382 ( .A1(n20002), .A2(n26130), .B1(n10628), .B2(n10081), .ZN(
        n20547) );
  NOR4_X2 U383 ( .A1(n10629), .A2(n10630), .A3(n10631), .A4(n10632), .ZN(
        n10628) );
  NAND4_X2 U384 ( .A1(n10633), .A2(n10634), .A3(n10635), .A4(n10636), .ZN(
        n10632) );
  AOI221_X2 U385 ( .B1(n10090), .B2(n25316), .C1(n10092), .C2(n24937), .A(
        n10639), .ZN(n10636) );
  OAI22_X2 U386 ( .A1(n19988), .A2(n10095), .B1(n19987), .B2(n10096), .ZN(
        n10639) );
  AOI221_X2 U389 ( .B1(n10097), .B2(n25315), .C1(n10099), .C2(n24936), .A(
        n10642), .ZN(n10635) );
  OAI22_X2 U390 ( .A1(n19994), .A2(n10102), .B1(n19993), .B2(n10103), .ZN(
        n10642) );
  AOI221_X2 U393 ( .B1(n10104), .B2(n25314), .C1(n10106), .C2(n24935), .A(
        n10645), .ZN(n10634) );
  OAI22_X2 U394 ( .A1(n19996), .A2(n10109), .B1(n19995), .B2(n10110), .ZN(
        n10645) );
  AOI221_X2 U397 ( .B1(n10111), .B2(n25313), .C1(n19945), .C2(n26139), .A(
        n10647), .ZN(n10633) );
  OAI22_X2 U398 ( .A1(n20000), .A2(n10115), .B1(n19999), .B2(n10116), .ZN(
        n10647) );
  NAND4_X2 U400 ( .A1(n10648), .A2(n10649), .A3(n10650), .A4(n10651), .ZN(
        n10631) );
  AOI221_X2 U401 ( .B1(n10121), .B2(n25355), .C1(n10123), .C2(n24934), .A(
        n10654), .ZN(n10651) );
  OAI22_X2 U402 ( .A1(n19972), .A2(n10126), .B1(n19971), .B2(n10127), .ZN(
        n10654) );
  AOI221_X2 U405 ( .B1(n10128), .B2(n28625), .C1(n10130), .C2(n28465), .A(
        n10657), .ZN(n10650) );
  OAI22_X2 U406 ( .A1(n19978), .A2(n10133), .B1(n19977), .B2(n10134), .ZN(
        n10657) );
  AOI221_X2 U409 ( .B1(n10135), .B2(n25312), .C1(n10137), .C2(n24933), .A(
        n10660), .ZN(n10649) );
  OAI22_X2 U410 ( .A1(n19980), .A2(n10140), .B1(n19979), .B2(n10141), .ZN(
        n10660) );
  AOI221_X2 U413 ( .B1(n10142), .B2(n25073), .C1(n10144), .C2(n25579), .A(
        n10663), .ZN(n10648) );
  OAI22_X2 U414 ( .A1(n19986), .A2(n10147), .B1(n19985), .B2(n10148), .ZN(
        n10663) );
  NAND4_X2 U417 ( .A1(n10664), .A2(n10665), .A3(n10666), .A4(n10667), .ZN(
        n10630) );
  AOI221_X2 U418 ( .B1(n19951), .B2(n10153), .C1(n19950), .C2(n10154), .A(
        n10668), .ZN(n10667) );
  OAI22_X2 U419 ( .A1(n10156), .A2(n28616), .B1(n10158), .B2(n28615), .ZN(
        n10668) );
  AOI221_X2 U420 ( .B1(n19947), .B2(n10160), .C1(n19946), .C2(n10161), .A(
        n10671), .ZN(n10666) );
  OAI22_X2 U421 ( .A1(n10163), .A2(n28323), .B1(n10165), .B2(n28322), .ZN(
        n10671) );
  AOI221_X2 U422 ( .B1(n19942), .B2(n10167), .C1(n19941), .C2(n10168), .A(
        n10674), .ZN(n10665) );
  OAI22_X2 U423 ( .A1(n10170), .A2(n28463), .B1(n10172), .B2(n28619), .ZN(
        n10674) );
  AOI221_X2 U424 ( .B1(n19938), .B2(n10174), .C1(n10175), .C2(n25578), .A(
        n10678), .ZN(n10664) );
  OAI22_X2 U425 ( .A1(n10178), .A2(n28203), .B1(n10180), .B2(n28202), .ZN(
        n10678) );
  NAND4_X2 U427 ( .A1(n10681), .A2(n10682), .A3(n10683), .A4(n10684), .ZN(
        n10629) );
  AOI221_X2 U428 ( .B1(n19969), .B2(n10186), .C1(n19968), .C2(n10187), .A(
        n10685), .ZN(n10684) );
  OAI22_X2 U429 ( .A1(n10189), .A2(n28623), .B1(n10191), .B2(n28621), .ZN(
        n10685) );
  AOI221_X2 U430 ( .B1(n19963), .B2(n10193), .C1(n19962), .C2(n10194), .A(
        n10688), .ZN(n10683) );
  OAI22_X2 U431 ( .A1(n10196), .A2(n28326), .B1(n10198), .B2(n28328), .ZN(
        n10688) );
  AOI221_X2 U432 ( .B1(n19959), .B2(n10200), .C1(n19958), .C2(n10201), .A(
        n10691), .ZN(n10682) );
  OAI22_X2 U433 ( .A1(n10203), .A2(n28460), .B1(n10205), .B2(n28459), .ZN(
        n10691) );
  AOI221_X2 U434 ( .B1(n19955), .B2(n10207), .C1(n19954), .C2(n10208), .A(
        n10694), .ZN(n10681) );
  OAI22_X2 U435 ( .A1(n10210), .A2(n28199), .B1(n10212), .B2(n28198), .ZN(
        n10694) );
  OAI22_X2 U436 ( .A1(n20067), .A2(n26130), .B1(n10697), .B2(n10081), .ZN(
        n20548) );
  NOR4_X2 U437 ( .A1(n10698), .A2(n10699), .A3(n10700), .A4(n10701), .ZN(
        n10697) );
  NAND4_X2 U438 ( .A1(n10702), .A2(n10703), .A3(n10704), .A4(n10705), .ZN(
        n10701) );
  AOI221_X2 U439 ( .B1(n10090), .B2(n25311), .C1(n10092), .C2(n24932), .A(
        n10708), .ZN(n10705) );
  OAI22_X2 U440 ( .A1(n20053), .A2(n10095), .B1(n20052), .B2(n10096), .ZN(
        n10708) );
  AOI221_X2 U443 ( .B1(n10097), .B2(n25310), .C1(n10099), .C2(n24931), .A(
        n10711), .ZN(n10704) );
  OAI22_X2 U444 ( .A1(n20059), .A2(n10102), .B1(n20058), .B2(n10103), .ZN(
        n10711) );
  AOI221_X2 U447 ( .B1(n10104), .B2(n25309), .C1(n10106), .C2(n24930), .A(
        n10714), .ZN(n10703) );
  OAI22_X2 U448 ( .A1(n20061), .A2(n10109), .B1(n20060), .B2(n10110), .ZN(
        n10714) );
  AOI221_X2 U451 ( .B1(n10111), .B2(n25308), .C1(n20010), .C2(n26139), .A(
        n10716), .ZN(n10702) );
  OAI22_X2 U452 ( .A1(n20065), .A2(n10115), .B1(n20064), .B2(n10116), .ZN(
        n10716) );
  NAND4_X2 U454 ( .A1(n10717), .A2(n10718), .A3(n10719), .A4(n10720), .ZN(
        n10700) );
  AOI221_X2 U455 ( .B1(n10121), .B2(n25354), .C1(n10123), .C2(n24929), .A(
        n10723), .ZN(n10720) );
  OAI22_X2 U456 ( .A1(n20037), .A2(n10126), .B1(n20036), .B2(n10127), .ZN(
        n10723) );
  AOI221_X2 U459 ( .B1(n10128), .B2(n28614), .C1(n10130), .C2(n28458), .A(
        n10726), .ZN(n10719) );
  OAI22_X2 U460 ( .A1(n20043), .A2(n10133), .B1(n20042), .B2(n10134), .ZN(
        n10726) );
  AOI221_X2 U463 ( .B1(n10135), .B2(n25307), .C1(n10137), .C2(n24928), .A(
        n10729), .ZN(n10718) );
  OAI22_X2 U464 ( .A1(n20045), .A2(n10140), .B1(n20044), .B2(n10141), .ZN(
        n10729) );
  AOI221_X2 U467 ( .B1(n10142), .B2(n25072), .C1(n10144), .C2(n25577), .A(
        n10732), .ZN(n10717) );
  OAI22_X2 U468 ( .A1(n20051), .A2(n10147), .B1(n20050), .B2(n10148), .ZN(
        n10732) );
  NAND4_X2 U471 ( .A1(n10733), .A2(n10734), .A3(n10735), .A4(n10736), .ZN(
        n10699) );
  AOI221_X2 U472 ( .B1(n20016), .B2(n10153), .C1(n20015), .C2(n10154), .A(
        n10737), .ZN(n10736) );
  OAI22_X2 U473 ( .A1(n10156), .A2(n28605), .B1(n10158), .B2(n28604), .ZN(
        n10737) );
  AOI221_X2 U474 ( .B1(n20012), .B2(n10160), .C1(n20011), .C2(n10161), .A(
        n10740), .ZN(n10735) );
  OAI22_X2 U475 ( .A1(n10163), .A2(n28315), .B1(n10165), .B2(n28314), .ZN(
        n10740) );
  AOI221_X2 U476 ( .B1(n20007), .B2(n10167), .C1(n20006), .C2(n10168), .A(
        n10743), .ZN(n10734) );
  OAI22_X2 U477 ( .A1(n10170), .A2(n28456), .B1(n10172), .B2(n28608), .ZN(
        n10743) );
  AOI221_X2 U478 ( .B1(n20003), .B2(n10174), .C1(n10175), .C2(n25576), .A(
        n10747), .ZN(n10733) );
  OAI22_X2 U479 ( .A1(n10178), .A2(n28195), .B1(n10180), .B2(n28194), .ZN(
        n10747) );
  NAND4_X2 U481 ( .A1(n10750), .A2(n10751), .A3(n10752), .A4(n10753), .ZN(
        n10698) );
  AOI221_X2 U482 ( .B1(n20034), .B2(n10186), .C1(n20033), .C2(n10187), .A(
        n10754), .ZN(n10753) );
  OAI22_X2 U483 ( .A1(n10189), .A2(n28612), .B1(n10191), .B2(n28610), .ZN(
        n10754) );
  AOI221_X2 U484 ( .B1(n20028), .B2(n10193), .C1(n20027), .C2(n10194), .A(
        n10757), .ZN(n10752) );
  OAI22_X2 U485 ( .A1(n10196), .A2(n28318), .B1(n10198), .B2(n28320), .ZN(
        n10757) );
  AOI221_X2 U486 ( .B1(n20024), .B2(n10200), .C1(n20023), .C2(n10201), .A(
        n10760), .ZN(n10751) );
  OAI22_X2 U487 ( .A1(n10203), .A2(n28453), .B1(n10205), .B2(n28452), .ZN(
        n10760) );
  AOI221_X2 U488 ( .B1(n20020), .B2(n10207), .C1(n20019), .C2(n10208), .A(
        n10763), .ZN(n10750) );
  OAI22_X2 U489 ( .A1(n10210), .A2(n28191), .B1(n10212), .B2(n28190), .ZN(
        n10763) );
  OAI22_X2 U490 ( .A1(n20132), .A2(n26130), .B1(n10766), .B2(n10081), .ZN(
        n20549) );
  NOR4_X2 U491 ( .A1(n10767), .A2(n10768), .A3(n10769), .A4(n10770), .ZN(
        n10766) );
  NAND4_X2 U492 ( .A1(n10771), .A2(n10772), .A3(n10773), .A4(n10774), .ZN(
        n10770) );
  AOI221_X2 U493 ( .B1(n10090), .B2(n25306), .C1(n10092), .C2(n24927), .A(
        n10777), .ZN(n10774) );
  OAI22_X2 U494 ( .A1(n20118), .A2(n10095), .B1(n20117), .B2(n10096), .ZN(
        n10777) );
  AOI221_X2 U497 ( .B1(n10097), .B2(n25305), .C1(n10099), .C2(n24926), .A(
        n10780), .ZN(n10773) );
  OAI22_X2 U498 ( .A1(n20124), .A2(n10102), .B1(n20123), .B2(n10103), .ZN(
        n10780) );
  AOI221_X2 U501 ( .B1(n10104), .B2(n25304), .C1(n10106), .C2(n24925), .A(
        n10783), .ZN(n10772) );
  OAI22_X2 U502 ( .A1(n20126), .A2(n10109), .B1(n20125), .B2(n10110), .ZN(
        n10783) );
  AOI221_X2 U505 ( .B1(n10111), .B2(n25303), .C1(n20075), .C2(n26139), .A(
        n10785), .ZN(n10771) );
  OAI22_X2 U506 ( .A1(n20130), .A2(n10115), .B1(n20129), .B2(n10116), .ZN(
        n10785) );
  NAND4_X2 U508 ( .A1(n10786), .A2(n10787), .A3(n10788), .A4(n10789), .ZN(
        n10769) );
  AOI221_X2 U509 ( .B1(n10121), .B2(n25353), .C1(n10123), .C2(n24924), .A(
        n10792), .ZN(n10789) );
  OAI22_X2 U510 ( .A1(n20102), .A2(n10126), .B1(n20101), .B2(n10127), .ZN(
        n10792) );
  AOI221_X2 U513 ( .B1(n10128), .B2(n28603), .C1(n10130), .C2(n28451), .A(
        n10795), .ZN(n10788) );
  OAI22_X2 U514 ( .A1(n20108), .A2(n10133), .B1(n20107), .B2(n10134), .ZN(
        n10795) );
  AOI221_X2 U517 ( .B1(n10135), .B2(n25302), .C1(n10137), .C2(n24923), .A(
        n10798), .ZN(n10787) );
  OAI22_X2 U518 ( .A1(n20110), .A2(n10140), .B1(n20109), .B2(n10141), .ZN(
        n10798) );
  AOI221_X2 U521 ( .B1(n10142), .B2(n25071), .C1(n10144), .C2(n25575), .A(
        n10801), .ZN(n10786) );
  OAI22_X2 U522 ( .A1(n20116), .A2(n10147), .B1(n20115), .B2(n10148), .ZN(
        n10801) );
  NAND4_X2 U525 ( .A1(n10802), .A2(n10803), .A3(n10804), .A4(n10805), .ZN(
        n10768) );
  AOI221_X2 U526 ( .B1(n20081), .B2(n10153), .C1(n20080), .C2(n10154), .A(
        n10806), .ZN(n10805) );
  OAI22_X2 U527 ( .A1(n10156), .A2(n28594), .B1(n10158), .B2(n28593), .ZN(
        n10806) );
  AOI221_X2 U528 ( .B1(n20077), .B2(n10160), .C1(n20076), .C2(n10161), .A(
        n10809), .ZN(n10804) );
  OAI22_X2 U529 ( .A1(n10163), .A2(n28307), .B1(n10165), .B2(n28306), .ZN(
        n10809) );
  AOI221_X2 U530 ( .B1(n20072), .B2(n10167), .C1(n20071), .C2(n10168), .A(
        n10812), .ZN(n10803) );
  OAI22_X2 U531 ( .A1(n10170), .A2(n28449), .B1(n10172), .B2(n28597), .ZN(
        n10812) );
  AOI221_X2 U532 ( .B1(n20068), .B2(n10174), .C1(n10175), .C2(n25574), .A(
        n10816), .ZN(n10802) );
  OAI22_X2 U533 ( .A1(n10178), .A2(n28187), .B1(n10180), .B2(n28186), .ZN(
        n10816) );
  NAND4_X2 U535 ( .A1(n10819), .A2(n10820), .A3(n10821), .A4(n10822), .ZN(
        n10767) );
  AOI221_X2 U536 ( .B1(n20099), .B2(n10186), .C1(n20098), .C2(n10187), .A(
        n10823), .ZN(n10822) );
  OAI22_X2 U537 ( .A1(n10189), .A2(n28601), .B1(n10191), .B2(n28599), .ZN(
        n10823) );
  AOI221_X2 U538 ( .B1(n20093), .B2(n10193), .C1(n20092), .C2(n10194), .A(
        n10826), .ZN(n10821) );
  OAI22_X2 U539 ( .A1(n10196), .A2(n28310), .B1(n10198), .B2(n28312), .ZN(
        n10826) );
  AOI221_X2 U540 ( .B1(n20089), .B2(n10200), .C1(n20088), .C2(n10201), .A(
        n10829), .ZN(n10820) );
  OAI22_X2 U541 ( .A1(n10203), .A2(n28446), .B1(n10205), .B2(n28445), .ZN(
        n10829) );
  AOI221_X2 U542 ( .B1(n20085), .B2(n10207), .C1(n20084), .C2(n10208), .A(
        n10832), .ZN(n10819) );
  OAI22_X2 U543 ( .A1(n10210), .A2(n28183), .B1(n10212), .B2(n28182), .ZN(
        n10832) );
  NAND4_X2 U546 ( .A1(n10840), .A2(n10841), .A3(n10842), .A4(n10843), .ZN(
        n10839) );
  AOI221_X2 U547 ( .B1(n10090), .B2(n25301), .C1(n10092), .C2(n24922), .A(
        n10846), .ZN(n10843) );
  OAI22_X2 U548 ( .A1(n20183), .A2(n10095), .B1(n20182), .B2(n10096), .ZN(
        n10846) );
  AOI221_X2 U551 ( .B1(n10097), .B2(n25300), .C1(n10099), .C2(n24921), .A(
        n10849), .ZN(n10842) );
  OAI22_X2 U552 ( .A1(n20189), .A2(n10102), .B1(n20188), .B2(n10103), .ZN(
        n10849) );
  AOI221_X2 U555 ( .B1(n10104), .B2(n25299), .C1(n10106), .C2(n24920), .A(
        n10852), .ZN(n10841) );
  OAI22_X2 U556 ( .A1(n20191), .A2(n10109), .B1(n20190), .B2(n10110), .ZN(
        n10852) );
  AOI221_X2 U559 ( .B1(n10111), .B2(n25298), .C1(n20140), .C2(n26139), .A(
        n10854), .ZN(n10840) );
  OAI22_X2 U560 ( .A1(n20195), .A2(n10115), .B1(n20194), .B2(n10116), .ZN(
        n10854) );
  NAND4_X2 U562 ( .A1(n10855), .A2(n10856), .A3(n10857), .A4(n10858), .ZN(
        n10838) );
  AOI221_X2 U563 ( .B1(n10121), .B2(n25352), .C1(n10123), .C2(n24919), .A(
        n10861), .ZN(n10858) );
  OAI22_X2 U564 ( .A1(n20167), .A2(n10126), .B1(n20166), .B2(n10127), .ZN(
        n10861) );
  AOI221_X2 U567 ( .B1(n10128), .B2(n28592), .C1(n10130), .C2(n28444), .A(
        n10864), .ZN(n10857) );
  OAI22_X2 U568 ( .A1(n20173), .A2(n10133), .B1(n20172), .B2(n10134), .ZN(
        n10864) );
  AOI221_X2 U571 ( .B1(n10135), .B2(n25297), .C1(n10137), .C2(n24918), .A(
        n10867), .ZN(n10856) );
  OAI22_X2 U572 ( .A1(n20175), .A2(n10140), .B1(n20174), .B2(n10141), .ZN(
        n10867) );
  AOI221_X2 U575 ( .B1(n10142), .B2(n25296), .C1(n10144), .C2(n24917), .A(
        n10870), .ZN(n10855) );
  OAI22_X2 U576 ( .A1(n20181), .A2(n10147), .B1(n20180), .B2(n10148), .ZN(
        n10870) );
  NAND4_X2 U579 ( .A1(n10871), .A2(n10872), .A3(n10873), .A4(n10874), .ZN(
        n10837) );
  AOI221_X2 U580 ( .B1(n20146), .B2(n10153), .C1(n20145), .C2(n10154), .A(
        n10875), .ZN(n10874) );
  OAI22_X2 U581 ( .A1(n10156), .A2(n28583), .B1(n10158), .B2(n28582), .ZN(
        n10875) );
  AOI221_X2 U582 ( .B1(n20142), .B2(n10160), .C1(n20141), .C2(n10161), .A(
        n10878), .ZN(n10873) );
  OAI22_X2 U583 ( .A1(n10163), .A2(n28299), .B1(n10165), .B2(n28298), .ZN(
        n10878) );
  AOI221_X2 U584 ( .B1(n20137), .B2(n10167), .C1(n20136), .C2(n10168), .A(
        n10881), .ZN(n10872) );
  OAI22_X2 U585 ( .A1(n10170), .A2(n28442), .B1(n10172), .B2(n28586), .ZN(
        n10881) );
  AOI221_X2 U586 ( .B1(n20133), .B2(n10174), .C1(n10175), .C2(n25264), .A(
        n10885), .ZN(n10871) );
  OAI22_X2 U587 ( .A1(n10178), .A2(n28179), .B1(n10180), .B2(n28178), .ZN(
        n10885) );
  NAND4_X2 U589 ( .A1(n10888), .A2(n10889), .A3(n10890), .A4(n10891), .ZN(
        n10836) );
  AOI221_X2 U590 ( .B1(n20164), .B2(n10186), .C1(n20163), .C2(n10187), .A(
        n10892), .ZN(n10891) );
  OAI22_X2 U591 ( .A1(n10189), .A2(n28590), .B1(n10191), .B2(n28588), .ZN(
        n10892) );
  AOI221_X2 U592 ( .B1(n20158), .B2(n10193), .C1(n20157), .C2(n10194), .A(
        n10895), .ZN(n10890) );
  OAI22_X2 U593 ( .A1(n10196), .A2(n28302), .B1(n10198), .B2(n28304), .ZN(
        n10895) );
  AOI221_X2 U594 ( .B1(n20154), .B2(n10200), .C1(n20153), .C2(n10201), .A(
        n10898), .ZN(n10889) );
  OAI22_X2 U595 ( .A1(n10203), .A2(n28439), .B1(n10205), .B2(n28438), .ZN(
        n10898) );
  AOI221_X2 U596 ( .B1(n20150), .B2(n10207), .C1(n20149), .C2(n10208), .A(
        n10901), .ZN(n10888) );
  OAI22_X2 U597 ( .A1(n10210), .A2(n28175), .B1(n10212), .B2(n28174), .ZN(
        n10901) );
  NAND4_X2 U600 ( .A1(n10909), .A2(n10910), .A3(n10911), .A4(n10912), .ZN(
        n10908) );
  AOI221_X2 U601 ( .B1(n10090), .B2(n25295), .C1(n10092), .C2(n24916), .A(
        n10915), .ZN(n10912) );
  OAI22_X2 U602 ( .A1(n20248), .A2(n10095), .B1(n20247), .B2(n10096), .ZN(
        n10915) );
  AOI221_X2 U605 ( .B1(n10097), .B2(n25294), .C1(n10099), .C2(n24915), .A(
        n10918), .ZN(n10911) );
  OAI22_X2 U606 ( .A1(n20254), .A2(n10102), .B1(n20253), .B2(n10103), .ZN(
        n10918) );
  AOI221_X2 U609 ( .B1(n10104), .B2(n25293), .C1(n10106), .C2(n24914), .A(
        n10921), .ZN(n10910) );
  OAI22_X2 U610 ( .A1(n20256), .A2(n10109), .B1(n20255), .B2(n10110), .ZN(
        n10921) );
  AOI221_X2 U613 ( .B1(n10111), .B2(n25292), .C1(n20205), .C2(n26139), .A(
        n10923), .ZN(n10909) );
  OAI22_X2 U614 ( .A1(n20260), .A2(n10115), .B1(n20259), .B2(n10116), .ZN(
        n10923) );
  NAND4_X2 U616 ( .A1(n10924), .A2(n10925), .A3(n10926), .A4(n10927), .ZN(
        n10907) );
  AOI221_X2 U617 ( .B1(n10121), .B2(n25351), .C1(n10123), .C2(n24913), .A(
        n10930), .ZN(n10927) );
  OAI22_X2 U618 ( .A1(n20232), .A2(n10126), .B1(n20231), .B2(n10127), .ZN(
        n10930) );
  AOI221_X2 U621 ( .B1(n10128), .B2(n28581), .C1(n10130), .C2(n28437), .A(
        n10933), .ZN(n10926) );
  OAI22_X2 U622 ( .A1(n20238), .A2(n10133), .B1(n20237), .B2(n10134), .ZN(
        n10933) );
  AOI221_X2 U625 ( .B1(n10135), .B2(n25291), .C1(n10137), .C2(n24912), .A(
        n10936), .ZN(n10925) );
  OAI22_X2 U626 ( .A1(n20240), .A2(n10140), .B1(n20239), .B2(n10141), .ZN(
        n10936) );
  AOI221_X2 U629 ( .B1(n10142), .B2(n25290), .C1(n10144), .C2(n24911), .A(
        n10939), .ZN(n10924) );
  OAI22_X2 U630 ( .A1(n20246), .A2(n10147), .B1(n20245), .B2(n10148), .ZN(
        n10939) );
  NAND4_X2 U633 ( .A1(n10940), .A2(n10941), .A3(n10942), .A4(n10943), .ZN(
        n10906) );
  AOI221_X2 U634 ( .B1(n20211), .B2(n10153), .C1(n20210), .C2(n10154), .A(
        n10944), .ZN(n10943) );
  OAI22_X2 U635 ( .A1(n10156), .A2(n28572), .B1(n10158), .B2(n28571), .ZN(
        n10944) );
  AOI221_X2 U636 ( .B1(n20207), .B2(n10160), .C1(n20206), .C2(n10161), .A(
        n10947), .ZN(n10942) );
  OAI22_X2 U637 ( .A1(n10163), .A2(n28291), .B1(n10165), .B2(n28290), .ZN(
        n10947) );
  AOI221_X2 U638 ( .B1(n20202), .B2(n10167), .C1(n20201), .C2(n10168), .A(
        n10950), .ZN(n10941) );
  OAI22_X2 U639 ( .A1(n10170), .A2(n28435), .B1(n10172), .B2(n28575), .ZN(
        n10950) );
  AOI221_X2 U640 ( .B1(n20198), .B2(n10174), .C1(n10175), .C2(n25573), .A(
        n10954), .ZN(n10940) );
  OAI22_X2 U641 ( .A1(n10178), .A2(n28171), .B1(n10180), .B2(n28170), .ZN(
        n10954) );
  NAND4_X2 U643 ( .A1(n10957), .A2(n10958), .A3(n10959), .A4(n10960), .ZN(
        n10905) );
  AOI221_X2 U644 ( .B1(n20229), .B2(n10186), .C1(n20228), .C2(n10187), .A(
        n10961), .ZN(n10960) );
  OAI22_X2 U645 ( .A1(n10189), .A2(n28579), .B1(n10191), .B2(n28577), .ZN(
        n10961) );
  AOI221_X2 U646 ( .B1(n20223), .B2(n10193), .C1(n20222), .C2(n10194), .A(
        n10964), .ZN(n10959) );
  OAI22_X2 U647 ( .A1(n10196), .A2(n28294), .B1(n10198), .B2(n28296), .ZN(
        n10964) );
  AOI221_X2 U648 ( .B1(n20219), .B2(n10200), .C1(n20218), .C2(n10201), .A(
        n10967), .ZN(n10958) );
  OAI22_X2 U649 ( .A1(n10203), .A2(n28432), .B1(n10205), .B2(n28431), .ZN(
        n10967) );
  AOI221_X2 U650 ( .B1(n20215), .B2(n10207), .C1(n20214), .C2(n10208), .A(
        n10970), .ZN(n10957) );
  OAI22_X2 U651 ( .A1(n10210), .A2(n28167), .B1(n10212), .B2(n28166), .ZN(
        n10970) );
  NAND4_X2 U654 ( .A1(n10978), .A2(n10979), .A3(n10980), .A4(n10981), .ZN(
        n10977) );
  AOI221_X2 U655 ( .B1(n10090), .B2(n25289), .C1(n10092), .C2(n28568), .A(
        n10984), .ZN(n10981) );
  OAI22_X2 U656 ( .A1(n20313), .A2(n10095), .B1(n20312), .B2(n10096), .ZN(
        n10984) );
  AOI221_X2 U659 ( .B1(n10097), .B2(n28567), .C1(n10099), .C2(n28566), .A(
        n10987), .ZN(n10980) );
  OAI22_X2 U660 ( .A1(n20319), .A2(n10102), .B1(n20318), .B2(n10103), .ZN(
        n10987) );
  AOI221_X2 U663 ( .B1(n10104), .B2(n25288), .C1(n10106), .C2(n28430), .A(
        n10990), .ZN(n10979) );
  OAI22_X2 U664 ( .A1(n20321), .A2(n10109), .B1(n20320), .B2(n10110), .ZN(
        n10990) );
  AOI221_X2 U667 ( .B1(n10111), .B2(n28429), .C1(n20270), .C2(n26139), .A(
        n10992), .ZN(n10978) );
  OAI22_X2 U668 ( .A1(n20325), .A2(n10115), .B1(n20324), .B2(n10116), .ZN(
        n10992) );
  NAND4_X2 U670 ( .A1(n10993), .A2(n10994), .A3(n10995), .A4(n10996), .ZN(
        n10976) );
  AOI221_X2 U671 ( .B1(n10121), .B2(n25350), .C1(n10123), .C2(n28570), .A(
        n10999), .ZN(n10996) );
  OAI22_X2 U672 ( .A1(n20297), .A2(n10126), .B1(n20296), .B2(n10127), .ZN(
        n10999) );
  AOI221_X2 U675 ( .B1(n10128), .B2(n28569), .C1(n10130), .C2(n28428), .A(
        n11002), .ZN(n10995) );
  OAI22_X2 U676 ( .A1(n20303), .A2(n10133), .B1(n20302), .B2(n10134), .ZN(
        n11002) );
  AOI221_X2 U679 ( .B1(n10135), .B2(n25287), .C1(n10137), .C2(n28427), .A(
        n11005), .ZN(n10994) );
  OAI22_X2 U680 ( .A1(n20305), .A2(n10140), .B1(n20304), .B2(n10141), .ZN(
        n11005) );
  AOI221_X2 U683 ( .B1(n10142), .B2(n28426), .C1(n10144), .C2(n28425), .A(
        n11008), .ZN(n10993) );
  OAI22_X2 U684 ( .A1(n20311), .A2(n10147), .B1(n20310), .B2(n10148), .ZN(
        n11008) );
  NAND4_X2 U687 ( .A1(n11009), .A2(n11010), .A3(n11011), .A4(n11012), .ZN(
        n10975) );
  AOI221_X2 U688 ( .B1(n20276), .B2(n10153), .C1(n20275), .C2(n10154), .A(
        n11013), .ZN(n11012) );
  OAI22_X2 U689 ( .A1(n10156), .A2(n28557), .B1(n10158), .B2(n28556), .ZN(
        n11013) );
  AOI221_X2 U690 ( .B1(n20272), .B2(n10160), .C1(n20271), .C2(n10161), .A(
        n11016), .ZN(n11011) );
  OAI22_X2 U691 ( .A1(n10163), .A2(n28283), .B1(n10165), .B2(n28282), .ZN(
        n11016) );
  AOI221_X2 U692 ( .B1(n20267), .B2(n10167), .C1(n20266), .C2(n10168), .A(
        n11019), .ZN(n11010) );
  OAI22_X2 U693 ( .A1(n10170), .A2(n28423), .B1(n10172), .B2(n28560), .ZN(
        n11019) );
  AOI221_X2 U694 ( .B1(n20263), .B2(n10174), .C1(n10175), .C2(n25572), .A(
        n11023), .ZN(n11009) );
  OAI22_X2 U695 ( .A1(n10178), .A2(n28163), .B1(n10180), .B2(n28162), .ZN(
        n11023) );
  NAND4_X2 U697 ( .A1(n11026), .A2(n11027), .A3(n11028), .A4(n11029), .ZN(
        n10974) );
  AOI221_X2 U698 ( .B1(n20294), .B2(n10186), .C1(n20293), .C2(n10187), .A(
        n11030), .ZN(n11029) );
  OAI22_X2 U699 ( .A1(n10189), .A2(n28564), .B1(n10191), .B2(n28562), .ZN(
        n11030) );
  AOI221_X2 U700 ( .B1(n20288), .B2(n10193), .C1(n20287), .C2(n10194), .A(
        n11033), .ZN(n11028) );
  OAI22_X2 U701 ( .A1(n10196), .A2(n28286), .B1(n10198), .B2(n28288), .ZN(
        n11033) );
  AOI221_X2 U702 ( .B1(n20284), .B2(n10200), .C1(n20283), .C2(n10201), .A(
        n11036), .ZN(n11027) );
  OAI22_X2 U703 ( .A1(n10203), .A2(n28420), .B1(n10205), .B2(n28419), .ZN(
        n11036) );
  AOI221_X2 U704 ( .B1(n20280), .B2(n10207), .C1(n20279), .C2(n10208), .A(
        n11039), .ZN(n11026) );
  OAI22_X2 U705 ( .A1(n10210), .A2(n28159), .B1(n10212), .B2(n28158), .ZN(
        n11039) );
  NAND4_X2 U708 ( .A1(n11047), .A2(n11048), .A3(n11049), .A4(n11050), .ZN(
        n11046) );
  AOI221_X2 U709 ( .B1(n10090), .B2(n25286), .C1(n10092), .C2(n28553), .A(
        n11053), .ZN(n11050) );
  OAI22_X2 U710 ( .A1(n20378), .A2(n10095), .B1(n20377), .B2(n10096), .ZN(
        n11053) );
  AOI221_X2 U713 ( .B1(n10097), .B2(n28552), .C1(n10099), .C2(n28551), .A(
        n11056), .ZN(n11049) );
  OAI22_X2 U714 ( .A1(n20384), .A2(n10102), .B1(n20383), .B2(n10103), .ZN(
        n11056) );
  AOI221_X2 U717 ( .B1(n10104), .B2(n25285), .C1(n10106), .C2(n28418), .A(
        n11059), .ZN(n11048) );
  OAI22_X2 U718 ( .A1(n20386), .A2(n10109), .B1(n20385), .B2(n10110), .ZN(
        n11059) );
  AOI221_X2 U721 ( .B1(n10111), .B2(n28417), .C1(n20335), .C2(n26139), .A(
        n11061), .ZN(n11047) );
  OAI22_X2 U722 ( .A1(n20390), .A2(n10115), .B1(n20389), .B2(n10116), .ZN(
        n11061) );
  NAND4_X2 U724 ( .A1(n11062), .A2(n11063), .A3(n11064), .A4(n11065), .ZN(
        n11045) );
  AOI221_X2 U725 ( .B1(n10121), .B2(n25349), .C1(n10123), .C2(n28555), .A(
        n11068), .ZN(n11065) );
  OAI22_X2 U726 ( .A1(n20362), .A2(n10126), .B1(n20361), .B2(n10127), .ZN(
        n11068) );
  AOI221_X2 U729 ( .B1(n10128), .B2(n28554), .C1(n10130), .C2(n28416), .A(
        n11071), .ZN(n11064) );
  OAI22_X2 U730 ( .A1(n20368), .A2(n10133), .B1(n20367), .B2(n10134), .ZN(
        n11071) );
  AOI221_X2 U733 ( .B1(n10135), .B2(n25284), .C1(n10137), .C2(n28415), .A(
        n11074), .ZN(n11063) );
  OAI22_X2 U734 ( .A1(n20370), .A2(n10140), .B1(n20369), .B2(n10141), .ZN(
        n11074) );
  AOI221_X2 U737 ( .B1(n10142), .B2(n28414), .C1(n10144), .C2(n28413), .A(
        n11077), .ZN(n11062) );
  OAI22_X2 U738 ( .A1(n20376), .A2(n10147), .B1(n20375), .B2(n10148), .ZN(
        n11077) );
  NAND4_X2 U741 ( .A1(n11078), .A2(n11079), .A3(n11080), .A4(n11081), .ZN(
        n11044) );
  AOI221_X2 U742 ( .B1(n20341), .B2(n10153), .C1(n20340), .C2(n10154), .A(
        n11082), .ZN(n11081) );
  OAI22_X2 U743 ( .A1(n10156), .A2(n28542), .B1(n10158), .B2(n28541), .ZN(
        n11082) );
  AOI221_X2 U744 ( .B1(n20337), .B2(n10160), .C1(n20336), .C2(n10161), .A(
        n11085), .ZN(n11080) );
  OAI22_X2 U745 ( .A1(n10163), .A2(n28275), .B1(n10165), .B2(n28274), .ZN(
        n11085) );
  AOI221_X2 U746 ( .B1(n20332), .B2(n10167), .C1(n20331), .C2(n10168), .A(
        n11088), .ZN(n11079) );
  OAI22_X2 U747 ( .A1(n10170), .A2(n28411), .B1(n10172), .B2(n28545), .ZN(
        n11088) );
  AOI221_X2 U748 ( .B1(n20328), .B2(n10174), .C1(n10175), .C2(n25571), .A(
        n11092), .ZN(n11078) );
  OAI22_X2 U749 ( .A1(n10178), .A2(n28155), .B1(n10180), .B2(n28154), .ZN(
        n11092) );
  NAND4_X2 U751 ( .A1(n11095), .A2(n11096), .A3(n11097), .A4(n11098), .ZN(
        n11043) );
  AOI221_X2 U752 ( .B1(n20359), .B2(n10186), .C1(n20358), .C2(n10187), .A(
        n11099), .ZN(n11098) );
  OAI22_X2 U753 ( .A1(n10189), .A2(n28549), .B1(n10191), .B2(n28547), .ZN(
        n11099) );
  AOI221_X2 U754 ( .B1(n20353), .B2(n10193), .C1(n20352), .C2(n10194), .A(
        n11102), .ZN(n11097) );
  OAI22_X2 U755 ( .A1(n10196), .A2(n28278), .B1(n10198), .B2(n28280), .ZN(
        n11102) );
  AOI221_X2 U756 ( .B1(n20349), .B2(n10200), .C1(n20348), .C2(n10201), .A(
        n11105), .ZN(n11096) );
  OAI22_X2 U757 ( .A1(n10203), .A2(n28408), .B1(n10205), .B2(n28407), .ZN(
        n11105) );
  AOI221_X2 U758 ( .B1(n20345), .B2(n10207), .C1(n20344), .C2(n10208), .A(
        n11108), .ZN(n11095) );
  OAI22_X2 U759 ( .A1(n10210), .A2(n28151), .B1(n10212), .B2(n28150), .ZN(
        n11108) );
  NAND4_X2 U762 ( .A1(n11116), .A2(n11117), .A3(n11118), .A4(n11119), .ZN(
        n11115) );
  AOI221_X2 U763 ( .B1(n10090), .B2(n25283), .C1(n10092), .C2(n28538), .A(
        n11122), .ZN(n11119) );
  OAI22_X2 U764 ( .A1(n20443), .A2(n10095), .B1(n20442), .B2(n10096), .ZN(
        n11122) );
  AOI221_X2 U767 ( .B1(n10097), .B2(n28537), .C1(n10099), .C2(n28536), .A(
        n11125), .ZN(n11118) );
  OAI22_X2 U768 ( .A1(n20449), .A2(n10102), .B1(n20448), .B2(n10103), .ZN(
        n11125) );
  AOI221_X2 U771 ( .B1(n10104), .B2(n25282), .C1(n10106), .C2(n28406), .A(
        n11128), .ZN(n11117) );
  OAI22_X2 U772 ( .A1(n20451), .A2(n10109), .B1(n20450), .B2(n10110), .ZN(
        n11128) );
  AOI221_X2 U775 ( .B1(n10111), .B2(n28405), .C1(n20400), .C2(n26139), .A(
        n11130), .ZN(n11116) );
  OAI22_X2 U776 ( .A1(n20455), .A2(n10115), .B1(n20454), .B2(n10116), .ZN(
        n11130) );
  NAND4_X2 U778 ( .A1(n11131), .A2(n11132), .A3(n11133), .A4(n11134), .ZN(
        n11114) );
  AOI221_X2 U779 ( .B1(n10121), .B2(n25348), .C1(n10123), .C2(n28540), .A(
        n11137), .ZN(n11134) );
  OAI22_X2 U780 ( .A1(n20427), .A2(n10126), .B1(n20426), .B2(n10127), .ZN(
        n11137) );
  AOI221_X2 U783 ( .B1(n10128), .B2(n28539), .C1(n10130), .C2(n28404), .A(
        n11140), .ZN(n11133) );
  OAI22_X2 U784 ( .A1(n20433), .A2(n10133), .B1(n20432), .B2(n10134), .ZN(
        n11140) );
  AOI221_X2 U787 ( .B1(n10135), .B2(n25281), .C1(n10137), .C2(n28403), .A(
        n11143), .ZN(n11132) );
  OAI22_X2 U788 ( .A1(n20435), .A2(n10140), .B1(n20434), .B2(n10141), .ZN(
        n11143) );
  AOI221_X2 U791 ( .B1(n10142), .B2(n28402), .C1(n10144), .C2(n28401), .A(
        n11146), .ZN(n11131) );
  OAI22_X2 U792 ( .A1(n20441), .A2(n10147), .B1(n20440), .B2(n10148), .ZN(
        n11146) );
  NAND4_X2 U795 ( .A1(n11147), .A2(n11148), .A3(n11149), .A4(n11150), .ZN(
        n11113) );
  AOI221_X2 U796 ( .B1(n20406), .B2(n10153), .C1(n20405), .C2(n10154), .A(
        n11151), .ZN(n11150) );
  OAI22_X2 U797 ( .A1(n10156), .A2(n28527), .B1(n10158), .B2(n28526), .ZN(
        n11151) );
  AOI221_X2 U798 ( .B1(n20402), .B2(n10160), .C1(n20401), .C2(n10161), .A(
        n11154), .ZN(n11149) );
  OAI22_X2 U799 ( .A1(n10163), .A2(n28267), .B1(n10165), .B2(n28266), .ZN(
        n11154) );
  AOI221_X2 U800 ( .B1(n20397), .B2(n10167), .C1(n20396), .C2(n10168), .A(
        n11157), .ZN(n11148) );
  OAI22_X2 U801 ( .A1(n10170), .A2(n28399), .B1(n10172), .B2(n28530), .ZN(
        n11157) );
  AOI221_X2 U802 ( .B1(n20393), .B2(n10174), .C1(n10175), .C2(n25263), .A(
        n11161), .ZN(n11147) );
  OAI22_X2 U803 ( .A1(n10178), .A2(n28147), .B1(n10180), .B2(n28146), .ZN(
        n11161) );
  NAND4_X2 U805 ( .A1(n11164), .A2(n11165), .A3(n11166), .A4(n11167), .ZN(
        n11112) );
  AOI221_X2 U806 ( .B1(n20424), .B2(n10186), .C1(n20423), .C2(n10187), .A(
        n11168), .ZN(n11167) );
  OAI22_X2 U807 ( .A1(n10189), .A2(n28534), .B1(n10191), .B2(n28532), .ZN(
        n11168) );
  AOI221_X2 U808 ( .B1(n20418), .B2(n10193), .C1(n20417), .C2(n10194), .A(
        n11171), .ZN(n11166) );
  OAI22_X2 U809 ( .A1(n10196), .A2(n28270), .B1(n10198), .B2(n28272), .ZN(
        n11171) );
  AOI221_X2 U810 ( .B1(n20414), .B2(n10200), .C1(n20413), .C2(n10201), .A(
        n11174), .ZN(n11165) );
  OAI22_X2 U811 ( .A1(n10203), .A2(n28396), .B1(n10205), .B2(n28395), .ZN(
        n11174) );
  AOI221_X2 U812 ( .B1(n20410), .B2(n10207), .C1(n20409), .C2(n10208), .A(
        n11177), .ZN(n11164) );
  OAI22_X2 U813 ( .A1(n10210), .A2(n28143), .B1(n10212), .B2(n28142), .ZN(
        n11177) );
  NAND4_X2 U816 ( .A1(n11185), .A2(n11186), .A3(n11187), .A4(n11188), .ZN(
        n11184) );
  AOI221_X2 U817 ( .B1(n10090), .B2(n25280), .C1(n10092), .C2(n28523), .A(
        n11191), .ZN(n11188) );
  OAI22_X2 U818 ( .A1(n20509), .A2(n10095), .B1(n20508), .B2(n10096), .ZN(
        n11191) );
  AOI221_X2 U825 ( .B1(n10097), .B2(n28522), .C1(n10099), .C2(n28521), .A(
        n11199), .ZN(n11187) );
  OAI22_X2 U826 ( .A1(n20515), .A2(n10102), .B1(n20514), .B2(n10103), .ZN(
        n11199) );
  AOI221_X2 U834 ( .B1(n10104), .B2(n25279), .C1(n10106), .C2(n28394), .A(
        n11206), .ZN(n11186) );
  OAI22_X2 U835 ( .A1(n20517), .A2(n10109), .B1(n20516), .B2(n10110), .ZN(
        n11206) );
  AOI221_X2 U842 ( .B1(n10111), .B2(n28393), .C1(n20466), .C2(n26139), .A(
        n11209), .ZN(n11185) );
  OAI22_X2 U843 ( .A1(n20521), .A2(n10115), .B1(n20520), .B2(n10116), .ZN(
        n11209) );
  NAND4_X2 U850 ( .A1(n11213), .A2(n11214), .A3(n11215), .A4(n11216), .ZN(
        n11183) );
  AOI221_X2 U851 ( .B1(n10121), .B2(n25347), .C1(n10123), .C2(n28525), .A(
        n11219), .ZN(n11216) );
  OAI22_X2 U852 ( .A1(n20493), .A2(n10126), .B1(n20492), .B2(n10127), .ZN(
        n11219) );
  AOI221_X2 U859 ( .B1(n10128), .B2(n28524), .C1(n10130), .C2(n28392), .A(
        n11224), .ZN(n11215) );
  OAI22_X2 U860 ( .A1(n20499), .A2(n10133), .B1(n20498), .B2(n10134), .ZN(
        n11224) );
  AOI221_X2 U867 ( .B1(n10135), .B2(n25278), .C1(n10137), .C2(n28391), .A(
        n11230), .ZN(n11214) );
  OAI22_X2 U868 ( .A1(n20501), .A2(n10140), .B1(n20500), .B2(n10141), .ZN(
        n11230) );
  AOI221_X2 U875 ( .B1(n10142), .B2(n28390), .C1(n10144), .C2(n28389), .A(
        n11234), .ZN(n11213) );
  OAI22_X2 U876 ( .A1(n20507), .A2(n10147), .B1(n20506), .B2(n10148), .ZN(
        n11234) );
  NAND4_X2 U886 ( .A1(n11237), .A2(n11238), .A3(n11239), .A4(n11240), .ZN(
        n11182) );
  AOI221_X2 U887 ( .B1(n20472), .B2(n10153), .C1(n20471), .C2(n10154), .A(
        n11241), .ZN(n11240) );
  OAI22_X2 U888 ( .A1(n10156), .A2(n28512), .B1(n10158), .B2(n28511), .ZN(
        n11241) );
  AOI221_X2 U893 ( .B1(n20468), .B2(n10160), .C1(n20467), .C2(n10161), .A(
        n11246), .ZN(n11239) );
  OAI22_X2 U894 ( .A1(n10163), .A2(n28259), .B1(n10165), .B2(n28258), .ZN(
        n11246) );
  NOR2_X2 U901 ( .A1(add_283_A_4_), .A2(n22414), .ZN(n11236) );
  AOI221_X2 U902 ( .B1(n20463), .B2(n10167), .C1(n20462), .C2(n10168), .A(
        n11250), .ZN(n11238) );
  OAI22_X2 U903 ( .A1(n10170), .A2(n28387), .B1(n10172), .B2(n28515), .ZN(
        n11250) );
  AOI221_X2 U908 ( .B1(n20459), .B2(n10174), .C1(n10175), .C2(n25570), .A(
        n11254), .ZN(n11237) );
  OAI22_X2 U909 ( .A1(n10178), .A2(n28139), .B1(n10180), .B2(n28138), .ZN(
        n11254) );
  NAND4_X2 U918 ( .A1(n11258), .A2(n11259), .A3(n11260), .A4(n11261), .ZN(
        n11181) );
  AOI221_X2 U919 ( .B1(n20490), .B2(n10186), .C1(n20489), .C2(n10187), .A(
        n11262), .ZN(n11261) );
  OAI22_X2 U920 ( .A1(n10189), .A2(n28519), .B1(n10191), .B2(n28517), .ZN(
        n11262) );
  AOI221_X2 U925 ( .B1(n20484), .B2(n10193), .C1(n20483), .C2(n10194), .A(
        n11267), .ZN(n11260) );
  OAI22_X2 U926 ( .A1(n10196), .A2(n28262), .B1(n10198), .B2(n28264), .ZN(
        n11267) );
  NOR2_X2 U931 ( .A1(add_283_A_0_), .A2(n22418), .ZN(n11235) );
  AOI221_X2 U935 ( .B1(n20480), .B2(n10200), .C1(n20479), .C2(n10201), .A(
        n11272), .ZN(n11259) );
  OAI22_X2 U936 ( .A1(n10203), .A2(n28384), .B1(n10205), .B2(n28383), .ZN(
        n11272) );
  AOI221_X2 U942 ( .B1(n20476), .B2(n10207), .C1(n20475), .C2(n10208), .A(
        n11278), .ZN(n11258) );
  OAI22_X2 U943 ( .A1(n10210), .A2(n28135), .B1(n10212), .B2(n28134), .ZN(
        n11278) );
  NOR2_X2 U953 ( .A1(add_283_A_1_), .A2(n22419), .ZN(n11212) );
  NOR2_X2 U954 ( .A1(add_283_A_5_), .A2(n22415), .ZN(n11202) );
  OAI22_X2 U960 ( .A1(n11283), .A2(n26279), .B1(n20528), .B2(n25959), .ZN(
        n20560) );
  OAI22_X2 U961 ( .A1(n11283), .A2(n26278), .B1(n20529), .B2(n25959), .ZN(
        n20561) );
  OAI22_X2 U962 ( .A1(n11283), .A2(n26277), .B1(n20530), .B2(n25959), .ZN(
        n20562) );
  OAI22_X2 U963 ( .A1(n11283), .A2(n26276), .B1(n20531), .B2(n25959), .ZN(
        n20563) );
  OAI22_X2 U964 ( .A1(n25958), .A2(n26275), .B1(n20532), .B2(n25959), .ZN(
        n20564) );
  OAI22_X2 U965 ( .A1(n25958), .A2(n26274), .B1(n20533), .B2(n25959), .ZN(
        n20565) );
  OAI22_X2 U966 ( .A1(n25958), .A2(n26273), .B1(n20534), .B2(n25959), .ZN(
        n20566) );
  OAI22_X2 U967 ( .A1(n25958), .A2(n26272), .B1(n20535), .B2(n25959), .ZN(
        n20567) );
  OAI22_X2 U968 ( .A1(n25958), .A2(n26271), .B1(n20536), .B2(n25959), .ZN(
        n20568) );
  OAI22_X2 U969 ( .A1(n25958), .A2(n26270), .B1(n20537), .B2(n25959), .ZN(
        n20569) );
  OAI22_X2 U970 ( .A1(n25958), .A2(n26269), .B1(n20538), .B2(n25959), .ZN(
        n20570) );
  OAI22_X2 U971 ( .A1(n25958), .A2(n26268), .B1(n20539), .B2(n25959), .ZN(
        n20571) );
  OAI22_X2 U973 ( .A1(n24846), .A2(n26220), .B1(n20432), .B2(n25956), .ZN(
        n20573) );
  OAI22_X2 U974 ( .A1(n25955), .A2(n26219), .B1(n20367), .B2(n25956), .ZN(
        n20574) );
  OAI22_X2 U975 ( .A1(n25955), .A2(n26218), .B1(n20302), .B2(n25956), .ZN(
        n20575) );
  OAI22_X2 U976 ( .A1(n24846), .A2(n26217), .B1(n20237), .B2(n25956), .ZN(
        n20576) );
  OAI22_X2 U977 ( .A1(n24846), .A2(n26216), .B1(n20172), .B2(n25956), .ZN(
        n20577) );
  OAI22_X2 U978 ( .A1(n24846), .A2(n26215), .B1(n20107), .B2(n25956), .ZN(
        n20578) );
  OAI22_X2 U979 ( .A1(n24846), .A2(n26214), .B1(n20042), .B2(n25956), .ZN(
        n20579) );
  OAI22_X2 U980 ( .A1(n24846), .A2(n26213), .B1(n19977), .B2(n25956), .ZN(
        n20580) );
  OAI22_X2 U981 ( .A1(n24846), .A2(n26212), .B1(n19912), .B2(n25956), .ZN(
        n20581) );
  OAI22_X2 U982 ( .A1(n24846), .A2(n26211), .B1(n19847), .B2(n25956), .ZN(
        n20582) );
  OAI22_X2 U983 ( .A1(n24846), .A2(n26210), .B1(n19782), .B2(n25956), .ZN(
        n20583) );
  OAI22_X2 U984 ( .A1(n25955), .A2(n26209), .B1(n19717), .B2(n25956), .ZN(
        n20584) );
  OAI22_X2 U985 ( .A1(n25955), .A2(n26208), .B1(n19652), .B2(n25956), .ZN(
        n20585) );
  OAI22_X2 U986 ( .A1(n25955), .A2(n26207), .B1(n19587), .B2(n25956), .ZN(
        n20586) );
  OAI22_X2 U988 ( .A1(n25955), .A2(n26206), .B1(n20494), .B2(n25956), .ZN(
        n20588) );
  OAI22_X2 U989 ( .A1(n25955), .A2(n26205), .B1(n20428), .B2(n25956), .ZN(
        n20589) );
  OAI22_X2 U990 ( .A1(n25955), .A2(n26204), .B1(n20363), .B2(n25956), .ZN(
        n20590) );
  OAI22_X2 U991 ( .A1(n25955), .A2(n26203), .B1(n20298), .B2(n25956), .ZN(
        n20591) );
  OAI22_X2 U992 ( .A1(n25955), .A2(n26202), .B1(n20233), .B2(n25956), .ZN(
        n20592) );
  OAI22_X2 U993 ( .A1(n25955), .A2(n26201), .B1(n20168), .B2(n25956), .ZN(
        n20593) );
  OAI22_X2 U994 ( .A1(n25955), .A2(n26200), .B1(n20103), .B2(n25956), .ZN(
        n20594) );
  OAI22_X2 U995 ( .A1(n25955), .A2(n26199), .B1(n20038), .B2(n25956), .ZN(
        n20595) );
  OAI22_X2 U996 ( .A1(n25955), .A2(n26198), .B1(n19973), .B2(n25956), .ZN(
        n20596) );
  OAI22_X2 U997 ( .A1(n25955), .A2(n26197), .B1(n19908), .B2(n25956), .ZN(
        n20597) );
  OAI22_X2 U998 ( .A1(n25955), .A2(n26196), .B1(n19843), .B2(n25956), .ZN(
        n20598) );
  OAI22_X2 U999 ( .A1(n25955), .A2(n26195), .B1(n19778), .B2(n25956), .ZN(
        n20599) );
  OAI22_X2 U1000 ( .A1(n25955), .A2(n26194), .B1(n19713), .B2(n25956), .ZN(
        n20600) );
  OAI22_X2 U1001 ( .A1(n24846), .A2(n26193), .B1(n19648), .B2(n25956), .ZN(
        n20601) );
  OAI22_X2 U1008 ( .A1(n20258), .A2(n25953), .B1(n26217), .B2(n25952), .ZN(
        n20608) );
  OAI22_X2 U1009 ( .A1(n20193), .A2(n25953), .B1(n26216), .B2(n25952), .ZN(
        n20609) );
  OAI22_X2 U1010 ( .A1(n20128), .A2(n25953), .B1(n26215), .B2(n25952), .ZN(
        n20610) );
  OAI22_X2 U1011 ( .A1(n20063), .A2(n25953), .B1(n26214), .B2(n25952), .ZN(
        n20611) );
  OAI22_X2 U1012 ( .A1(n19998), .A2(n25953), .B1(n26213), .B2(n25952), .ZN(
        n20612) );
  OAI22_X2 U1013 ( .A1(n19933), .A2(n25953), .B1(n26212), .B2(n25952), .ZN(
        n20613) );
  OAI22_X2 U1014 ( .A1(n19868), .A2(n25953), .B1(n26211), .B2(n24864), .ZN(
        n20614) );
  OAI22_X2 U1015 ( .A1(n19803), .A2(n25953), .B1(n26210), .B2(n24864), .ZN(
        n20615) );
  OAI22_X2 U1016 ( .A1(n19738), .A2(n25953), .B1(n26209), .B2(n25952), .ZN(
        n20616) );
  OAI22_X2 U1017 ( .A1(n19673), .A2(n25953), .B1(n26208), .B2(n25952), .ZN(
        n20617) );
  OAI22_X2 U1018 ( .A1(n19608), .A2(n25953), .B1(n26207), .B2(n25952), .ZN(
        n20618) );
  OAI22_X2 U1020 ( .A1(n20515), .A2(n25953), .B1(n25952), .B2(n26266), .ZN(
        n20620) );
  OAI22_X2 U1021 ( .A1(n20449), .A2(n25953), .B1(n25952), .B2(n26265), .ZN(
        n20621) );
  OAI22_X2 U1022 ( .A1(n20384), .A2(n25953), .B1(n24864), .B2(n26264), .ZN(
        n20622) );
  OAI22_X2 U1023 ( .A1(n20319), .A2(n25953), .B1(n24864), .B2(n26263), .ZN(
        n20623) );
  OAI22_X2 U1024 ( .A1(n20254), .A2(n25953), .B1(n24864), .B2(n26262), .ZN(
        n20624) );
  OAI22_X2 U1025 ( .A1(n20189), .A2(n25953), .B1(n25952), .B2(n26261), .ZN(
        n20625) );
  OAI22_X2 U1026 ( .A1(n20124), .A2(n25953), .B1(n24864), .B2(n26260), .ZN(
        n20626) );
  OAI22_X2 U1027 ( .A1(n20059), .A2(n25953), .B1(n24864), .B2(n26259), .ZN(
        n20627) );
  OAI22_X2 U1028 ( .A1(n19994), .A2(n25953), .B1(n24864), .B2(n26258), .ZN(
        n20628) );
  OAI22_X2 U1029 ( .A1(n19929), .A2(n25953), .B1(n24864), .B2(n26257), .ZN(
        n20629) );
  OAI22_X2 U1030 ( .A1(n19864), .A2(n25953), .B1(n24864), .B2(n26256), .ZN(
        n20630) );
  OAI22_X2 U1031 ( .A1(n19799), .A2(n25953), .B1(n25952), .B2(n26255), .ZN(
        n20631) );
  OAI22_X2 U1032 ( .A1(n19734), .A2(n25953), .B1(n25952), .B2(n26254), .ZN(
        n20632) );
  OAI22_X2 U1033 ( .A1(n19669), .A2(n25953), .B1(n25952), .B2(n26253), .ZN(
        n20633) );
  OAI22_X2 U1034 ( .A1(n19604), .A2(n25953), .B1(n25952), .B2(n26252), .ZN(
        n20634) );
  OAI22_X2 U1036 ( .A1(n20495), .A2(n25951), .B1(n24845), .B2(n26251), .ZN(
        n20636) );
  OAI22_X2 U1037 ( .A1(n20429), .A2(n25951), .B1(n24845), .B2(n26250), .ZN(
        n20637) );
  OAI22_X2 U1038 ( .A1(n20364), .A2(n25950), .B1(n24845), .B2(n26249), .ZN(
        n20638) );
  OAI22_X2 U1039 ( .A1(n20299), .A2(n25950), .B1(n24845), .B2(n26248), .ZN(
        n20639) );
  OAI22_X2 U1040 ( .A1(n20234), .A2(n25950), .B1(n25949), .B2(n26247), .ZN(
        n20640) );
  OAI22_X2 U1041 ( .A1(n20169), .A2(n25950), .B1(n25949), .B2(n26246), .ZN(
        n20641) );
  OAI22_X2 U1042 ( .A1(n20104), .A2(n25950), .B1(n25949), .B2(n26245), .ZN(
        n20642) );
  OAI22_X2 U1043 ( .A1(n20039), .A2(n25950), .B1(n25949), .B2(n26244), .ZN(
        n20643) );
  OAI22_X2 U1044 ( .A1(n19974), .A2(n25950), .B1(n24845), .B2(n26243), .ZN(
        n20644) );
  OAI22_X2 U1045 ( .A1(n19909), .A2(n25950), .B1(n25949), .B2(n26242), .ZN(
        n20645) );
  OAI22_X2 U1046 ( .A1(n19844), .A2(n25950), .B1(n25949), .B2(n26241), .ZN(
        n20646) );
  OAI22_X2 U1047 ( .A1(n19779), .A2(n25950), .B1(n25949), .B2(n26240), .ZN(
        n20647) );
  OAI22_X2 U1048 ( .A1(n19714), .A2(n25950), .B1(n25949), .B2(n26239), .ZN(
        n20648) );
  OAI22_X2 U1049 ( .A1(n19649), .A2(n25950), .B1(n25949), .B2(n26238), .ZN(
        n20649) );
  OAI22_X2 U1050 ( .A1(n19584), .A2(n25950), .B1(n25949), .B2(n26237), .ZN(
        n20650) );
  OAI22_X2 U1052 ( .A1(n20491), .A2(n25950), .B1(n26206), .B2(n25949), .ZN(
        n20652) );
  OAI22_X2 U1053 ( .A1(n20425), .A2(n25950), .B1(n26205), .B2(n25949), .ZN(
        n20653) );
  OAI22_X2 U1054 ( .A1(n20360), .A2(n25950), .B1(n26204), .B2(n25949), .ZN(
        n20654) );
  OAI22_X2 U1055 ( .A1(n20295), .A2(n25950), .B1(n26203), .B2(n25949), .ZN(
        n20655) );
  OAI22_X2 U1056 ( .A1(n20230), .A2(n25950), .B1(n26202), .B2(n25949), .ZN(
        n20656) );
  OAI22_X2 U1057 ( .A1(n20165), .A2(n25950), .B1(n26201), .B2(n25949), .ZN(
        n20657) );
  OAI22_X2 U1058 ( .A1(n20100), .A2(n25950), .B1(n26200), .B2(n25949), .ZN(
        n20658) );
  OAI22_X2 U1059 ( .A1(n20035), .A2(n25950), .B1(n26199), .B2(n25949), .ZN(
        n20659) );
  OAI22_X2 U1060 ( .A1(n19970), .A2(n25950), .B1(n26198), .B2(n25949), .ZN(
        n20660) );
  OAI22_X2 U1061 ( .A1(n19905), .A2(n25950), .B1(n26197), .B2(n25949), .ZN(
        n20661) );
  OAI22_X2 U1062 ( .A1(n19840), .A2(n25950), .B1(n26196), .B2(n25949), .ZN(
        n20662) );
  OAI22_X2 U1063 ( .A1(n19775), .A2(n25950), .B1(n26195), .B2(n25949), .ZN(
        n20663) );
  OAI22_X2 U1064 ( .A1(n19710), .A2(n25950), .B1(n26194), .B2(n24845), .ZN(
        n20664) );
  OAI22_X2 U1065 ( .A1(n19645), .A2(n25950), .B1(n26193), .B2(n25949), .ZN(
        n20665) );
  OAI22_X2 U1066 ( .A1(n19580), .A2(n25950), .B1(n26192), .B2(n24845), .ZN(
        n20666) );
  OAI22_X2 U1072 ( .A1(n20250), .A2(n25947), .B1(n26247), .B2(n25946), .ZN(
        n20672) );
  OAI22_X2 U1073 ( .A1(n20185), .A2(n25947), .B1(n26246), .B2(n25946), .ZN(
        n20673) );
  OAI22_X2 U1074 ( .A1(n20120), .A2(n25947), .B1(n26245), .B2(n24844), .ZN(
        n20674) );
  OAI22_X2 U1075 ( .A1(n20055), .A2(n25947), .B1(n26244), .B2(n24844), .ZN(
        n20675) );
  OAI22_X2 U1076 ( .A1(n19990), .A2(n25947), .B1(n26243), .B2(n24844), .ZN(
        n20676) );
  OAI22_X2 U1077 ( .A1(n19925), .A2(n25947), .B1(n26242), .B2(n24844), .ZN(
        n20677) );
  OAI22_X2 U1078 ( .A1(n19860), .A2(n25947), .B1(n26241), .B2(n24844), .ZN(
        n20678) );
  OAI22_X2 U1079 ( .A1(n19795), .A2(n25947), .B1(n26240), .B2(n24844), .ZN(
        n20679) );
  OAI22_X2 U1080 ( .A1(n19730), .A2(n25947), .B1(n26239), .B2(n25946), .ZN(
        n20680) );
  OAI22_X2 U1081 ( .A1(n19665), .A2(n25947), .B1(n26238), .B2(n25946), .ZN(
        n20681) );
  OAI22_X2 U1082 ( .A1(n19600), .A2(n25947), .B1(n26237), .B2(n25946), .ZN(
        n20682) );
  OAI22_X2 U1084 ( .A1(n20507), .A2(n25947), .B1(n26206), .B2(n25946), .ZN(
        n20684) );
  OAI22_X2 U1085 ( .A1(n20441), .A2(n25947), .B1(n26205), .B2(n25946), .ZN(
        n20685) );
  OAI22_X2 U1086 ( .A1(n20376), .A2(n25947), .B1(n26204), .B2(n24844), .ZN(
        n20686) );
  OAI22_X2 U1087 ( .A1(n20311), .A2(n25947), .B1(n26203), .B2(n24844), .ZN(
        n20687) );
  OAI22_X2 U1088 ( .A1(n20246), .A2(n25947), .B1(n26202), .B2(n24844), .ZN(
        n20688) );
  OAI22_X2 U1089 ( .A1(n20181), .A2(n25947), .B1(n26201), .B2(n24844), .ZN(
        n20689) );
  OAI22_X2 U1090 ( .A1(n20116), .A2(n25947), .B1(n26200), .B2(n24844), .ZN(
        n20690) );
  OAI22_X2 U1091 ( .A1(n20051), .A2(n25947), .B1(n26199), .B2(n25946), .ZN(
        n20691) );
  OAI22_X2 U1092 ( .A1(n19986), .A2(n25947), .B1(n26198), .B2(n25946), .ZN(
        n20692) );
  OAI22_X2 U1093 ( .A1(n19921), .A2(n25947), .B1(n26197), .B2(n25946), .ZN(
        n20693) );
  OAI22_X2 U1094 ( .A1(n19856), .A2(n25947), .B1(n26196), .B2(n25946), .ZN(
        n20694) );
  OAI22_X2 U1095 ( .A1(n19791), .A2(n25947), .B1(n26195), .B2(n25946), .ZN(
        n20695) );
  OAI22_X2 U1096 ( .A1(n19726), .A2(n25947), .B1(n26194), .B2(n25946), .ZN(
        n20696) );
  OAI22_X2 U1097 ( .A1(n19661), .A2(n25947), .B1(n26193), .B2(n24844), .ZN(
        n20697) );
  OAI22_X2 U1098 ( .A1(n19596), .A2(n25947), .B1(n26192), .B2(n24844), .ZN(
        n20698) );
  OAI22_X2 U1104 ( .A1(n20242), .A2(n25944), .B1(n26217), .B2(n25943), .ZN(
        n20704) );
  OAI22_X2 U1105 ( .A1(n20177), .A2(n25944), .B1(n26216), .B2(n25943), .ZN(
        n20705) );
  OAI22_X2 U1106 ( .A1(n20112), .A2(n25944), .B1(n26215), .B2(n25943), .ZN(
        n20706) );
  OAI22_X2 U1107 ( .A1(n20047), .A2(n25944), .B1(n26214), .B2(n24843), .ZN(
        n20707) );
  OAI22_X2 U1108 ( .A1(n19982), .A2(n25944), .B1(n26213), .B2(n24843), .ZN(
        n20708) );
  OAI22_X2 U1109 ( .A1(n19917), .A2(n25944), .B1(n26212), .B2(n24843), .ZN(
        n20709) );
  OAI22_X2 U1110 ( .A1(n19852), .A2(n25944), .B1(n26211), .B2(n24843), .ZN(
        n20710) );
  OAI22_X2 U1111 ( .A1(n19787), .A2(n25944), .B1(n26210), .B2(n24843), .ZN(
        n20711) );
  OAI22_X2 U1112 ( .A1(n19722), .A2(n25944), .B1(n26209), .B2(n25943), .ZN(
        n20712) );
  OAI22_X2 U1113 ( .A1(n19657), .A2(n25944), .B1(n26208), .B2(n25943), .ZN(
        n20713) );
  OAI22_X2 U1114 ( .A1(n19592), .A2(n25944), .B1(n26207), .B2(n25943), .ZN(
        n20714) );
  OAI22_X2 U1116 ( .A1(n20499), .A2(n25944), .B1(n26266), .B2(n24843), .ZN(
        n20716) );
  OAI22_X2 U1117 ( .A1(n20433), .A2(n25944), .B1(n26265), .B2(n24843), .ZN(
        n20717) );
  OAI22_X2 U1118 ( .A1(n20368), .A2(n25944), .B1(n26264), .B2(n24843), .ZN(
        n20718) );
  OAI22_X2 U1119 ( .A1(n20303), .A2(n25944), .B1(n26263), .B2(n24843), .ZN(
        n20719) );
  OAI22_X2 U1120 ( .A1(n20238), .A2(n25944), .B1(n26262), .B2(n24843), .ZN(
        n20720) );
  OAI22_X2 U1121 ( .A1(n20173), .A2(n25944), .B1(n26261), .B2(n25943), .ZN(
        n20721) );
  OAI22_X2 U1122 ( .A1(n20108), .A2(n25944), .B1(n26260), .B2(n25943), .ZN(
        n20722) );
  OAI22_X2 U1123 ( .A1(n20043), .A2(n25944), .B1(n26259), .B2(n25943), .ZN(
        n20723) );
  OAI22_X2 U1124 ( .A1(n19978), .A2(n25944), .B1(n26258), .B2(n25943), .ZN(
        n20724) );
  OAI22_X2 U1125 ( .A1(n19913), .A2(n25944), .B1(n26257), .B2(n25943), .ZN(
        n20725) );
  OAI22_X2 U1126 ( .A1(n19848), .A2(n25944), .B1(n26256), .B2(n25943), .ZN(
        n20726) );
  OAI22_X2 U1127 ( .A1(n19783), .A2(n25944), .B1(n26255), .B2(n24843), .ZN(
        n20727) );
  OAI22_X2 U1128 ( .A1(n19718), .A2(n25944), .B1(n26254), .B2(n25943), .ZN(
        n20728) );
  OAI22_X2 U1129 ( .A1(n19653), .A2(n25944), .B1(n26253), .B2(n24843), .ZN(
        n20729) );
  OAI22_X2 U1130 ( .A1(n19588), .A2(n25944), .B1(n26252), .B2(n24843), .ZN(
        n20730) );
  OAI22_X2 U1136 ( .A1(n20259), .A2(n25941), .B1(n26217), .B2(n25940), .ZN(
        n20736) );
  OAI22_X2 U1137 ( .A1(n20194), .A2(n25941), .B1(n26216), .B2(n25940), .ZN(
        n20737) );
  OAI22_X2 U1138 ( .A1(n20129), .A2(n25941), .B1(n26215), .B2(n25940), .ZN(
        n20738) );
  OAI22_X2 U1139 ( .A1(n20064), .A2(n25941), .B1(n26214), .B2(n24842), .ZN(
        n20739) );
  OAI22_X2 U1140 ( .A1(n19999), .A2(n25941), .B1(n26213), .B2(n24842), .ZN(
        n20740) );
  OAI22_X2 U1141 ( .A1(n19934), .A2(n25941), .B1(n26212), .B2(n24842), .ZN(
        n20741) );
  OAI22_X2 U1142 ( .A1(n19869), .A2(n25941), .B1(n26211), .B2(n24842), .ZN(
        n20742) );
  OAI22_X2 U1143 ( .A1(n19804), .A2(n25941), .B1(n26210), .B2(n24842), .ZN(
        n20743) );
  OAI22_X2 U1144 ( .A1(n19739), .A2(n25941), .B1(n26209), .B2(n25940), .ZN(
        n20744) );
  OAI22_X2 U1145 ( .A1(n19674), .A2(n25941), .B1(n26208), .B2(n24842), .ZN(
        n20745) );
  OAI22_X2 U1146 ( .A1(n19609), .A2(n25941), .B1(n26207), .B2(n24842), .ZN(
        n20746) );
  OAI22_X2 U1148 ( .A1(n20516), .A2(n25941), .B1(n26266), .B2(n24842), .ZN(
        n20748) );
  OAI22_X2 U1149 ( .A1(n20450), .A2(n25941), .B1(n26265), .B2(n24842), .ZN(
        n20749) );
  OAI22_X2 U1150 ( .A1(n20385), .A2(n25941), .B1(n26264), .B2(n24842), .ZN(
        n20750) );
  OAI22_X2 U1151 ( .A1(n20320), .A2(n25941), .B1(n26263), .B2(n25940), .ZN(
        n20751) );
  OAI22_X2 U1152 ( .A1(n20255), .A2(n25941), .B1(n26262), .B2(n25940), .ZN(
        n20752) );
  OAI22_X2 U1153 ( .A1(n20190), .A2(n25941), .B1(n26261), .B2(n25940), .ZN(
        n20753) );
  OAI22_X2 U1154 ( .A1(n20125), .A2(n25941), .B1(n26260), .B2(n25940), .ZN(
        n20754) );
  OAI22_X2 U1155 ( .A1(n20060), .A2(n25941), .B1(n26259), .B2(n25940), .ZN(
        n20755) );
  OAI22_X2 U1156 ( .A1(n19995), .A2(n25941), .B1(n26258), .B2(n25940), .ZN(
        n20756) );
  OAI22_X2 U1157 ( .A1(n19930), .A2(n25941), .B1(n26257), .B2(n25940), .ZN(
        n20757) );
  OAI22_X2 U1158 ( .A1(n19865), .A2(n25941), .B1(n26256), .B2(n25940), .ZN(
        n20758) );
  OAI22_X2 U1159 ( .A1(n19800), .A2(n25941), .B1(n26255), .B2(n24842), .ZN(
        n20759) );
  OAI22_X2 U1160 ( .A1(n19735), .A2(n25941), .B1(n26254), .B2(n25940), .ZN(
        n20760) );
  OAI22_X2 U1161 ( .A1(n19670), .A2(n25941), .B1(n26253), .B2(n24842), .ZN(
        n20761) );
  OAI22_X2 U1162 ( .A1(n19605), .A2(n25941), .B1(n26252), .B2(n24842), .ZN(
        n20762) );
  OAI22_X2 U1164 ( .A1(n20496), .A2(n25938), .B1(n26251), .B2(n25937), .ZN(
        n20764) );
  OAI22_X2 U1165 ( .A1(n20430), .A2(n25939), .B1(n26250), .B2(n25937), .ZN(
        n20765) );
  OAI22_X2 U1172 ( .A1(n19975), .A2(n25938), .B1(n26243), .B2(n24841), .ZN(
        n20772) );
  OAI22_X2 U1173 ( .A1(n19910), .A2(n25938), .B1(n26242), .B2(n24841), .ZN(
        n20773) );
  OAI22_X2 U1174 ( .A1(n19845), .A2(n25938), .B1(n26241), .B2(n24841), .ZN(
        n20774) );
  OAI22_X2 U1175 ( .A1(n19780), .A2(n25938), .B1(n26240), .B2(n24841), .ZN(
        n20775) );
  OAI22_X2 U1176 ( .A1(n19715), .A2(n25938), .B1(n26239), .B2(n25937), .ZN(
        n20776) );
  OAI22_X2 U1177 ( .A1(n19650), .A2(n25938), .B1(n26238), .B2(n25937), .ZN(
        n20777) );
  OAI22_X2 U1178 ( .A1(n19585), .A2(n25938), .B1(n26237), .B2(n25937), .ZN(
        n20778) );
  OAI22_X2 U1180 ( .A1(n20492), .A2(n25938), .B1(n26206), .B2(n24841), .ZN(
        n20780) );
  OAI22_X2 U1181 ( .A1(n20426), .A2(n25938), .B1(n26205), .B2(n24841), .ZN(
        n20781) );
  OAI22_X2 U1182 ( .A1(n20361), .A2(n25938), .B1(n26204), .B2(n24841), .ZN(
        n20782) );
  OAI22_X2 U1183 ( .A1(n20296), .A2(n25938), .B1(n26203), .B2(n24841), .ZN(
        n20783) );
  OAI22_X2 U1184 ( .A1(n20231), .A2(n25938), .B1(n26202), .B2(n24841), .ZN(
        n20784) );
  OAI22_X2 U1185 ( .A1(n20166), .A2(n25938), .B1(n26201), .B2(n25937), .ZN(
        n20785) );
  OAI22_X2 U1186 ( .A1(n20101), .A2(n25938), .B1(n26200), .B2(n25937), .ZN(
        n20786) );
  OAI22_X2 U1187 ( .A1(n20036), .A2(n25938), .B1(n26199), .B2(n25937), .ZN(
        n20787) );
  OAI22_X2 U1188 ( .A1(n19971), .A2(n25938), .B1(n26198), .B2(n25937), .ZN(
        n20788) );
  OAI22_X2 U1189 ( .A1(n19906), .A2(n25938), .B1(n26197), .B2(n25937), .ZN(
        n20789) );
  OAI22_X2 U1190 ( .A1(n19841), .A2(n25938), .B1(n26196), .B2(n25937), .ZN(
        n20790) );
  OAI22_X2 U1191 ( .A1(n19776), .A2(n25938), .B1(n26195), .B2(n25937), .ZN(
        n20791) );
  OAI22_X2 U1192 ( .A1(n19711), .A2(n25938), .B1(n26194), .B2(n25937), .ZN(
        n20792) );
  OAI22_X2 U1193 ( .A1(n19646), .A2(n25938), .B1(n26193), .B2(n24841), .ZN(
        n20793) );
  OAI22_X2 U1194 ( .A1(n19581), .A2(n25938), .B1(n26192), .B2(n24841), .ZN(
        n20794) );
  OAI22_X2 U1200 ( .A1(n20251), .A2(n25935), .B1(n26247), .B2(n25934), .ZN(
        n20800) );
  OAI22_X2 U1201 ( .A1(n20186), .A2(n25935), .B1(n26246), .B2(n25934), .ZN(
        n20801) );
  OAI22_X2 U1202 ( .A1(n20121), .A2(n25935), .B1(n26245), .B2(n24889), .ZN(
        n20802) );
  OAI22_X2 U1203 ( .A1(n20056), .A2(n25935), .B1(n26244), .B2(n24889), .ZN(
        n20803) );
  OAI22_X2 U1204 ( .A1(n19991), .A2(n25935), .B1(n26243), .B2(n24889), .ZN(
        n20804) );
  OAI22_X2 U1205 ( .A1(n19926), .A2(n25935), .B1(n26242), .B2(n24889), .ZN(
        n20805) );
  OAI22_X2 U1206 ( .A1(n19861), .A2(n25935), .B1(n26241), .B2(n24889), .ZN(
        n20806) );
  OAI22_X2 U1207 ( .A1(n19796), .A2(n25935), .B1(n26240), .B2(n24889), .ZN(
        n20807) );
  OAI22_X2 U1208 ( .A1(n19731), .A2(n25935), .B1(n26239), .B2(n25934), .ZN(
        n20808) );
  OAI22_X2 U1209 ( .A1(n19666), .A2(n25935), .B1(n26238), .B2(n25934), .ZN(
        n20809) );
  OAI22_X2 U1210 ( .A1(n19601), .A2(n25935), .B1(n26237), .B2(n25934), .ZN(
        n20810) );
  OAI22_X2 U1212 ( .A1(n20508), .A2(n25935), .B1(n26206), .B2(n24889), .ZN(
        n20812) );
  OAI22_X2 U1213 ( .A1(n20442), .A2(n25935), .B1(n26205), .B2(n24889), .ZN(
        n20813) );
  OAI22_X2 U1214 ( .A1(n20377), .A2(n25935), .B1(n26204), .B2(n24889), .ZN(
        n20814) );
  OAI22_X2 U1215 ( .A1(n20312), .A2(n25935), .B1(n26203), .B2(n24889), .ZN(
        n20815) );
  OAI22_X2 U1216 ( .A1(n20247), .A2(n25935), .B1(n26202), .B2(n24889), .ZN(
        n20816) );
  OAI22_X2 U1217 ( .A1(n20182), .A2(n25935), .B1(n26201), .B2(n25934), .ZN(
        n20817) );
  OAI22_X2 U1218 ( .A1(n20117), .A2(n25935), .B1(n26200), .B2(n25934), .ZN(
        n20818) );
  OAI22_X2 U1219 ( .A1(n20052), .A2(n25935), .B1(n26199), .B2(n25934), .ZN(
        n20819) );
  OAI22_X2 U1220 ( .A1(n19987), .A2(n25935), .B1(n26198), .B2(n25934), .ZN(
        n20820) );
  OAI22_X2 U1221 ( .A1(n19922), .A2(n25935), .B1(n26197), .B2(n25934), .ZN(
        n20821) );
  OAI22_X2 U1222 ( .A1(n19857), .A2(n25935), .B1(n26196), .B2(n25934), .ZN(
        n20822) );
  OAI22_X2 U1223 ( .A1(n19792), .A2(n25935), .B1(n26195), .B2(n25934), .ZN(
        n20823) );
  OAI22_X2 U1224 ( .A1(n19727), .A2(n25935), .B1(n26194), .B2(n25934), .ZN(
        n20824) );
  OAI22_X2 U1225 ( .A1(n19662), .A2(n25935), .B1(n26193), .B2(n24889), .ZN(
        n20825) );
  OAI22_X2 U1226 ( .A1(n19597), .A2(n25935), .B1(n26192), .B2(n24889), .ZN(
        n20826) );
  OAI22_X2 U1232 ( .A1(n20243), .A2(n25932), .B1(n26217), .B2(n25931), .ZN(
        n20832) );
  OAI22_X2 U1233 ( .A1(n20178), .A2(n25932), .B1(n26216), .B2(n25931), .ZN(
        n20833) );
  OAI22_X2 U1234 ( .A1(n20113), .A2(n25932), .B1(n26215), .B2(n25931), .ZN(
        n20834) );
  OAI22_X2 U1235 ( .A1(n20048), .A2(n25932), .B1(n26214), .B2(n24840), .ZN(
        n20835) );
  OAI22_X2 U1236 ( .A1(n19983), .A2(n25932), .B1(n26213), .B2(n24840), .ZN(
        n20836) );
  OAI22_X2 U1237 ( .A1(n19918), .A2(n25932), .B1(n26212), .B2(n24840), .ZN(
        n20837) );
  OAI22_X2 U1238 ( .A1(n19853), .A2(n25932), .B1(n26211), .B2(n24840), .ZN(
        n20838) );
  OAI22_X2 U1239 ( .A1(n19788), .A2(n25932), .B1(n26210), .B2(n24840), .ZN(
        n20839) );
  OAI22_X2 U1240 ( .A1(n19723), .A2(n25932), .B1(n26209), .B2(n25931), .ZN(
        n20840) );
  OAI22_X2 U1241 ( .A1(n19658), .A2(n25932), .B1(n26208), .B2(n24840), .ZN(
        n20841) );
  OAI22_X2 U1242 ( .A1(n19593), .A2(n25932), .B1(n26207), .B2(n24840), .ZN(
        n20842) );
  OAI22_X2 U1244 ( .A1(n20500), .A2(n25932), .B1(n26266), .B2(n24840), .ZN(
        n20844) );
  OAI22_X2 U1245 ( .A1(n20434), .A2(n25932), .B1(n26265), .B2(n24840), .ZN(
        n20845) );
  OAI22_X2 U1246 ( .A1(n20369), .A2(n25932), .B1(n26264), .B2(n24840), .ZN(
        n20846) );
  OAI22_X2 U1247 ( .A1(n20304), .A2(n25932), .B1(n26263), .B2(n25931), .ZN(
        n20847) );
  OAI22_X2 U1248 ( .A1(n20239), .A2(n25932), .B1(n26262), .B2(n25931), .ZN(
        n20848) );
  OAI22_X2 U1249 ( .A1(n20174), .A2(n25932), .B1(n26261), .B2(n25931), .ZN(
        n20849) );
  OAI22_X2 U1250 ( .A1(n20109), .A2(n25932), .B1(n26260), .B2(n25931), .ZN(
        n20850) );
  OAI22_X2 U1251 ( .A1(n20044), .A2(n25932), .B1(n26259), .B2(n25931), .ZN(
        n20851) );
  OAI22_X2 U1252 ( .A1(n19979), .A2(n25932), .B1(n26258), .B2(n25931), .ZN(
        n20852) );
  OAI22_X2 U1253 ( .A1(n19914), .A2(n25932), .B1(n26257), .B2(n25931), .ZN(
        n20853) );
  OAI22_X2 U1254 ( .A1(n19849), .A2(n25932), .B1(n26256), .B2(n25931), .ZN(
        n20854) );
  OAI22_X2 U1255 ( .A1(n19784), .A2(n25932), .B1(n26255), .B2(n24840), .ZN(
        n20855) );
  OAI22_X2 U1256 ( .A1(n19719), .A2(n25932), .B1(n26254), .B2(n25931), .ZN(
        n20856) );
  OAI22_X2 U1257 ( .A1(n19654), .A2(n25932), .B1(n26253), .B2(n24840), .ZN(
        n20857) );
  OAI22_X2 U1258 ( .A1(n19589), .A2(n25932), .B1(n26252), .B2(n24840), .ZN(
        n20858) );
  OAI22_X2 U1264 ( .A1(n20261), .A2(n25929), .B1(n26217), .B2(n25928), .ZN(
        n20864) );
  OAI22_X2 U1265 ( .A1(n20196), .A2(n25929), .B1(n26216), .B2(n25928), .ZN(
        n20865) );
  OAI22_X2 U1266 ( .A1(n20131), .A2(n25929), .B1(n26215), .B2(n25928), .ZN(
        n20866) );
  OAI22_X2 U1267 ( .A1(n20066), .A2(n25929), .B1(n26214), .B2(n24839), .ZN(
        n20867) );
  OAI22_X2 U1268 ( .A1(n20001), .A2(n25929), .B1(n26213), .B2(n24839), .ZN(
        n20868) );
  OAI22_X2 U1269 ( .A1(n19936), .A2(n25929), .B1(n26212), .B2(n24839), .ZN(
        n20869) );
  OAI22_X2 U1270 ( .A1(n19871), .A2(n25929), .B1(n26211), .B2(n24839), .ZN(
        n20870) );
  OAI22_X2 U1271 ( .A1(n19806), .A2(n25929), .B1(n26210), .B2(n24839), .ZN(
        n20871) );
  OAI22_X2 U1272 ( .A1(n19741), .A2(n25929), .B1(n26209), .B2(n25928), .ZN(
        n20872) );
  OAI22_X2 U1273 ( .A1(n19676), .A2(n25929), .B1(n26208), .B2(n25928), .ZN(
        n20873) );
  OAI22_X2 U1274 ( .A1(n19611), .A2(n25929), .B1(n26207), .B2(n25928), .ZN(
        n20874) );
  OAI22_X2 U1276 ( .A1(n20518), .A2(n25929), .B1(n26266), .B2(n24839), .ZN(
        n20876) );
  OAI22_X2 U1277 ( .A1(n20452), .A2(n25929), .B1(n26265), .B2(n24839), .ZN(
        n20877) );
  OAI22_X2 U1278 ( .A1(n20387), .A2(n25929), .B1(n26264), .B2(n24839), .ZN(
        n20878) );
  OAI22_X2 U1279 ( .A1(n20322), .A2(n25929), .B1(n26263), .B2(n24839), .ZN(
        n20879) );
  OAI22_X2 U1280 ( .A1(n20257), .A2(n25929), .B1(n26262), .B2(n24839), .ZN(
        n20880) );
  OAI22_X2 U1281 ( .A1(n20192), .A2(n25929), .B1(n26261), .B2(n25928), .ZN(
        n20881) );
  OAI22_X2 U1282 ( .A1(n20127), .A2(n25929), .B1(n26260), .B2(n25928), .ZN(
        n20882) );
  OAI22_X2 U1283 ( .A1(n20062), .A2(n25929), .B1(n26259), .B2(n25928), .ZN(
        n20883) );
  OAI22_X2 U1284 ( .A1(n19997), .A2(n25929), .B1(n26258), .B2(n25928), .ZN(
        n20884) );
  OAI22_X2 U1285 ( .A1(n19932), .A2(n25929), .B1(n26257), .B2(n25928), .ZN(
        n20885) );
  OAI22_X2 U1286 ( .A1(n19867), .A2(n25929), .B1(n26256), .B2(n25928), .ZN(
        n20886) );
  OAI22_X2 U1287 ( .A1(n19802), .A2(n25929), .B1(n26255), .B2(n24839), .ZN(
        n20887) );
  OAI22_X2 U1288 ( .A1(n19737), .A2(n25929), .B1(n26254), .B2(n25928), .ZN(
        n20888) );
  OAI22_X2 U1289 ( .A1(n19672), .A2(n25929), .B1(n26253), .B2(n24839), .ZN(
        n20889) );
  OAI22_X2 U1290 ( .A1(n19607), .A2(n25929), .B1(n26252), .B2(n24839), .ZN(
        n20890) );
  OAI22_X2 U1296 ( .A1(n20253), .A2(n25926), .B1(n26247), .B2(n25925), .ZN(
        n20896) );
  OAI22_X2 U1297 ( .A1(n20188), .A2(n25926), .B1(n26246), .B2(n25925), .ZN(
        n20897) );
  OAI22_X2 U1298 ( .A1(n20123), .A2(n25926), .B1(n26245), .B2(n24838), .ZN(
        n20898) );
  OAI22_X2 U1299 ( .A1(n20058), .A2(n25926), .B1(n26244), .B2(n24838), .ZN(
        n20899) );
  OAI22_X2 U1300 ( .A1(n19993), .A2(n25926), .B1(n26243), .B2(n24838), .ZN(
        n20900) );
  OAI22_X2 U1301 ( .A1(n19928), .A2(n25926), .B1(n26242), .B2(n24838), .ZN(
        n20901) );
  OAI22_X2 U1302 ( .A1(n19863), .A2(n25926), .B1(n26241), .B2(n24838), .ZN(
        n20902) );
  OAI22_X2 U1303 ( .A1(n19798), .A2(n25926), .B1(n26240), .B2(n24838), .ZN(
        n20903) );
  OAI22_X2 U1304 ( .A1(n19733), .A2(n25926), .B1(n26239), .B2(n25925), .ZN(
        n20904) );
  OAI22_X2 U1305 ( .A1(n19668), .A2(n25926), .B1(n26238), .B2(n25925), .ZN(
        n20905) );
  OAI22_X2 U1306 ( .A1(n19603), .A2(n25926), .B1(n26237), .B2(n25925), .ZN(
        n20906) );
  OAI22_X2 U1308 ( .A1(n20510), .A2(n25926), .B1(n26206), .B2(n25925), .ZN(
        n20908) );
  OAI22_X2 U1309 ( .A1(n20444), .A2(n25926), .B1(n26205), .B2(n25925), .ZN(
        n20909) );
  OAI22_X2 U1310 ( .A1(n20379), .A2(n25926), .B1(n26204), .B2(n24838), .ZN(
        n20910) );
  OAI22_X2 U1311 ( .A1(n20314), .A2(n25926), .B1(n26203), .B2(n24838), .ZN(
        n20911) );
  OAI22_X2 U1312 ( .A1(n20249), .A2(n25926), .B1(n26202), .B2(n24838), .ZN(
        n20912) );
  OAI22_X2 U1313 ( .A1(n20184), .A2(n25926), .B1(n26201), .B2(n24838), .ZN(
        n20913) );
  OAI22_X2 U1314 ( .A1(n20119), .A2(n25926), .B1(n26200), .B2(n24838), .ZN(
        n20914) );
  OAI22_X2 U1315 ( .A1(n20054), .A2(n25926), .B1(n26199), .B2(n25925), .ZN(
        n20915) );
  OAI22_X2 U1316 ( .A1(n19989), .A2(n25926), .B1(n26198), .B2(n25925), .ZN(
        n20916) );
  OAI22_X2 U1317 ( .A1(n19924), .A2(n25926), .B1(n26197), .B2(n25925), .ZN(
        n20917) );
  OAI22_X2 U1318 ( .A1(n19859), .A2(n25926), .B1(n26196), .B2(n25925), .ZN(
        n20918) );
  OAI22_X2 U1319 ( .A1(n19794), .A2(n25926), .B1(n26195), .B2(n25925), .ZN(
        n20919) );
  OAI22_X2 U1320 ( .A1(n19729), .A2(n25926), .B1(n26194), .B2(n25925), .ZN(
        n20920) );
  OAI22_X2 U1321 ( .A1(n19664), .A2(n25926), .B1(n26193), .B2(n24838), .ZN(
        n20921) );
  OAI22_X2 U1322 ( .A1(n19599), .A2(n25926), .B1(n26192), .B2(n24838), .ZN(
        n20922) );
  OAI22_X2 U1328 ( .A1(n20245), .A2(n25923), .B1(n26217), .B2(n25922), .ZN(
        n20928) );
  OAI22_X2 U1329 ( .A1(n20180), .A2(n25923), .B1(n26216), .B2(n25922), .ZN(
        n20929) );
  OAI22_X2 U1330 ( .A1(n20115), .A2(n25923), .B1(n26215), .B2(n25922), .ZN(
        n20930) );
  OAI22_X2 U1331 ( .A1(n20050), .A2(n25923), .B1(n26214), .B2(n24837), .ZN(
        n20931) );
  OAI22_X2 U1332 ( .A1(n19985), .A2(n25923), .B1(n26213), .B2(n24837), .ZN(
        n20932) );
  OAI22_X2 U1333 ( .A1(n19920), .A2(n25923), .B1(n26212), .B2(n24837), .ZN(
        n20933) );
  OAI22_X2 U1334 ( .A1(n19855), .A2(n25923), .B1(n26211), .B2(n24837), .ZN(
        n20934) );
  OAI22_X2 U1335 ( .A1(n19790), .A2(n25923), .B1(n26210), .B2(n24837), .ZN(
        n20935) );
  OAI22_X2 U1336 ( .A1(n19725), .A2(n25923), .B1(n26209), .B2(n25922), .ZN(
        n20936) );
  OAI22_X2 U1337 ( .A1(n19660), .A2(n25923), .B1(n26208), .B2(n25922), .ZN(
        n20937) );
  OAI22_X2 U1338 ( .A1(n19595), .A2(n25923), .B1(n26207), .B2(n25922), .ZN(
        n20938) );
  OAI22_X2 U1340 ( .A1(n20502), .A2(n25923), .B1(n26266), .B2(n24837), .ZN(
        n20940) );
  OAI22_X2 U1341 ( .A1(n20436), .A2(n25923), .B1(n26265), .B2(n24837), .ZN(
        n20941) );
  OAI22_X2 U1342 ( .A1(n20371), .A2(n25923), .B1(n26264), .B2(n24837), .ZN(
        n20942) );
  OAI22_X2 U1343 ( .A1(n20306), .A2(n25923), .B1(n26263), .B2(n24837), .ZN(
        n20943) );
  OAI22_X2 U1344 ( .A1(n20241), .A2(n25923), .B1(n26262), .B2(n24837), .ZN(
        n20944) );
  OAI22_X2 U1345 ( .A1(n20176), .A2(n25923), .B1(n26261), .B2(n25922), .ZN(
        n20945) );
  OAI22_X2 U1346 ( .A1(n20111), .A2(n25923), .B1(n26260), .B2(n25922), .ZN(
        n20946) );
  OAI22_X2 U1347 ( .A1(n20046), .A2(n25923), .B1(n26259), .B2(n25922), .ZN(
        n20947) );
  OAI22_X2 U1348 ( .A1(n19981), .A2(n25923), .B1(n26258), .B2(n25922), .ZN(
        n20948) );
  OAI22_X2 U1349 ( .A1(n19916), .A2(n25923), .B1(n26257), .B2(n25922), .ZN(
        n20949) );
  OAI22_X2 U1350 ( .A1(n19851), .A2(n25923), .B1(n26256), .B2(n25922), .ZN(
        n20950) );
  OAI22_X2 U1351 ( .A1(n19786), .A2(n25923), .B1(n26255), .B2(n24837), .ZN(
        n20951) );
  OAI22_X2 U1352 ( .A1(n19721), .A2(n25923), .B1(n26254), .B2(n25922), .ZN(
        n20952) );
  OAI22_X2 U1353 ( .A1(n19656), .A2(n25923), .B1(n26253), .B2(n24837), .ZN(
        n20953) );
  OAI22_X2 U1354 ( .A1(n19591), .A2(n25923), .B1(n26252), .B2(n24837), .ZN(
        n20954) );
  OAI22_X2 U1360 ( .A1(n20260), .A2(n25920), .B1(n26217), .B2(n25919), .ZN(
        n20960) );
  OAI22_X2 U1361 ( .A1(n20195), .A2(n25920), .B1(n26216), .B2(n25919), .ZN(
        n20961) );
  OAI22_X2 U1362 ( .A1(n20130), .A2(n25920), .B1(n26215), .B2(n25919), .ZN(
        n20962) );
  OAI22_X2 U1363 ( .A1(n20065), .A2(n25920), .B1(n26214), .B2(n24836), .ZN(
        n20963) );
  OAI22_X2 U1364 ( .A1(n20000), .A2(n25920), .B1(n26213), .B2(n24836), .ZN(
        n20964) );
  OAI22_X2 U1365 ( .A1(n19935), .A2(n25920), .B1(n26212), .B2(n24836), .ZN(
        n20965) );
  OAI22_X2 U1366 ( .A1(n19870), .A2(n25920), .B1(n26211), .B2(n24836), .ZN(
        n20966) );
  OAI22_X2 U1367 ( .A1(n19805), .A2(n25920), .B1(n26210), .B2(n24836), .ZN(
        n20967) );
  OAI22_X2 U1368 ( .A1(n19740), .A2(n25920), .B1(n26209), .B2(n25919), .ZN(
        n20968) );
  OAI22_X2 U1369 ( .A1(n19675), .A2(n25920), .B1(n26208), .B2(n24836), .ZN(
        n20969) );
  OAI22_X2 U1370 ( .A1(n19610), .A2(n25920), .B1(n26207), .B2(n24836), .ZN(
        n20970) );
  OAI22_X2 U1372 ( .A1(n20517), .A2(n25920), .B1(n26266), .B2(n24836), .ZN(
        n20972) );
  OAI22_X2 U1373 ( .A1(n20451), .A2(n25920), .B1(n26265), .B2(n24836), .ZN(
        n20973) );
  OAI22_X2 U1374 ( .A1(n20386), .A2(n25920), .B1(n26264), .B2(n24836), .ZN(
        n20974) );
  OAI22_X2 U1375 ( .A1(n20321), .A2(n25920), .B1(n26263), .B2(n25919), .ZN(
        n20975) );
  OAI22_X2 U1376 ( .A1(n20256), .A2(n25920), .B1(n26262), .B2(n25919), .ZN(
        n20976) );
  OAI22_X2 U1377 ( .A1(n20191), .A2(n25920), .B1(n26261), .B2(n25919), .ZN(
        n20977) );
  OAI22_X2 U1378 ( .A1(n20126), .A2(n25920), .B1(n26260), .B2(n25919), .ZN(
        n20978) );
  OAI22_X2 U1379 ( .A1(n20061), .A2(n25920), .B1(n26259), .B2(n25919), .ZN(
        n20979) );
  OAI22_X2 U1380 ( .A1(n19996), .A2(n25920), .B1(n26258), .B2(n25919), .ZN(
        n20980) );
  OAI22_X2 U1381 ( .A1(n19931), .A2(n25920), .B1(n26257), .B2(n25919), .ZN(
        n20981) );
  OAI22_X2 U1382 ( .A1(n19866), .A2(n25920), .B1(n26256), .B2(n25919), .ZN(
        n20982) );
  OAI22_X2 U1383 ( .A1(n19801), .A2(n25920), .B1(n26255), .B2(n24836), .ZN(
        n20983) );
  OAI22_X2 U1384 ( .A1(n19736), .A2(n25920), .B1(n26254), .B2(n25919), .ZN(
        n20984) );
  OAI22_X2 U1385 ( .A1(n19671), .A2(n25920), .B1(n26253), .B2(n24836), .ZN(
        n20985) );
  OAI22_X2 U1386 ( .A1(n19606), .A2(n25920), .B1(n26252), .B2(n24836), .ZN(
        n20986) );
  OAI22_X2 U1388 ( .A1(n20497), .A2(n25918), .B1(n26221), .B2(n25916), .ZN(
        n20988) );
  OAI22_X2 U1390 ( .A1(n20366), .A2(n25917), .B1(n26219), .B2(n25916), .ZN(
        n20990) );
  OAI22_X2 U1396 ( .A1(n19976), .A2(n25917), .B1(n26213), .B2(n24834), .ZN(
        n20996) );
  OAI22_X2 U1397 ( .A1(n19911), .A2(n25917), .B1(n26212), .B2(n24834), .ZN(
        n20997) );
  OAI22_X2 U1398 ( .A1(n19846), .A2(n25917), .B1(n26211), .B2(n24834), .ZN(
        n20998) );
  OAI22_X2 U1399 ( .A1(n19781), .A2(n25917), .B1(n26210), .B2(n24834), .ZN(
        n20999) );
  OAI22_X2 U1400 ( .A1(n19716), .A2(n25917), .B1(n26209), .B2(n24834), .ZN(
        n21000) );
  OAI22_X2 U1401 ( .A1(n19651), .A2(n25917), .B1(n26208), .B2(n25916), .ZN(
        n21001) );
  OAI22_X2 U1402 ( .A1(n19586), .A2(n25917), .B1(n26207), .B2(n25916), .ZN(
        n21002) );
  OAI22_X2 U1404 ( .A1(n20493), .A2(n25917), .B1(n26206), .B2(n25916), .ZN(
        n21004) );
  OAI22_X2 U1405 ( .A1(n20427), .A2(n25917), .B1(n26205), .B2(n25916), .ZN(
        n21005) );
  OAI22_X2 U1406 ( .A1(n20362), .A2(n25917), .B1(n26204), .B2(n25916), .ZN(
        n21006) );
  OAI22_X2 U1407 ( .A1(n20297), .A2(n25917), .B1(n26203), .B2(n24834), .ZN(
        n21007) );
  OAI22_X2 U1408 ( .A1(n20232), .A2(n25917), .B1(n26202), .B2(n24834), .ZN(
        n21008) );
  OAI22_X2 U1409 ( .A1(n20167), .A2(n25917), .B1(n26201), .B2(n24834), .ZN(
        n21009) );
  OAI22_X2 U1410 ( .A1(n20102), .A2(n25917), .B1(n26200), .B2(n24834), .ZN(
        n21010) );
  OAI22_X2 U1411 ( .A1(n20037), .A2(n25917), .B1(n26199), .B2(n25916), .ZN(
        n21011) );
  OAI22_X2 U1412 ( .A1(n19972), .A2(n25917), .B1(n26198), .B2(n25916), .ZN(
        n21012) );
  OAI22_X2 U1413 ( .A1(n19907), .A2(n25917), .B1(n26197), .B2(n25916), .ZN(
        n21013) );
  OAI22_X2 U1414 ( .A1(n19842), .A2(n25917), .B1(n26196), .B2(n25916), .ZN(
        n21014) );
  OAI22_X2 U1415 ( .A1(n19777), .A2(n25917), .B1(n26195), .B2(n25916), .ZN(
        n21015) );
  OAI22_X2 U1416 ( .A1(n19712), .A2(n25917), .B1(n26194), .B2(n25916), .ZN(
        n21016) );
  OAI22_X2 U1417 ( .A1(n19647), .A2(n25917), .B1(n26193), .B2(n25916), .ZN(
        n21017) );
  OAI22_X2 U1418 ( .A1(n19582), .A2(n25917), .B1(n26192), .B2(n25916), .ZN(
        n21018) );
  OAI22_X2 U1424 ( .A1(n20252), .A2(n25914), .B1(n26247), .B2(n25913), .ZN(
        n21024) );
  OAI22_X2 U1425 ( .A1(n20187), .A2(n25914), .B1(n26246), .B2(n25913), .ZN(
        n21025) );
  OAI22_X2 U1426 ( .A1(n20122), .A2(n25914), .B1(n26245), .B2(n24888), .ZN(
        n21026) );
  OAI22_X2 U1427 ( .A1(n20057), .A2(n25914), .B1(n26244), .B2(n24888), .ZN(
        n21027) );
  OAI22_X2 U1428 ( .A1(n19992), .A2(n25914), .B1(n26243), .B2(n24888), .ZN(
        n21028) );
  OAI22_X2 U1429 ( .A1(n19927), .A2(n25914), .B1(n26242), .B2(n24888), .ZN(
        n21029) );
  OAI22_X2 U1430 ( .A1(n19862), .A2(n25914), .B1(n26241), .B2(n24888), .ZN(
        n21030) );
  OAI22_X2 U1431 ( .A1(n19797), .A2(n25914), .B1(n26240), .B2(n24888), .ZN(
        n21031) );
  OAI22_X2 U1432 ( .A1(n19732), .A2(n25914), .B1(n26239), .B2(n25913), .ZN(
        n21032) );
  OAI22_X2 U1433 ( .A1(n19667), .A2(n25914), .B1(n26238), .B2(n25913), .ZN(
        n21033) );
  OAI22_X2 U1434 ( .A1(n19602), .A2(n25914), .B1(n26237), .B2(n25913), .ZN(
        n21034) );
  OAI22_X2 U1436 ( .A1(n20509), .A2(n25914), .B1(n26206), .B2(n24888), .ZN(
        n21036) );
  OAI22_X2 U1437 ( .A1(n20443), .A2(n25914), .B1(n26205), .B2(n24888), .ZN(
        n21037) );
  OAI22_X2 U1438 ( .A1(n20378), .A2(n25914), .B1(n26204), .B2(n24888), .ZN(
        n21038) );
  OAI22_X2 U1439 ( .A1(n20313), .A2(n25914), .B1(n26203), .B2(n24888), .ZN(
        n21039) );
  OAI22_X2 U1440 ( .A1(n20248), .A2(n25914), .B1(n26202), .B2(n24888), .ZN(
        n21040) );
  OAI22_X2 U1441 ( .A1(n20183), .A2(n25914), .B1(n26201), .B2(n25913), .ZN(
        n21041) );
  OAI22_X2 U1442 ( .A1(n20118), .A2(n25914), .B1(n26200), .B2(n25913), .ZN(
        n21042) );
  OAI22_X2 U1443 ( .A1(n20053), .A2(n25914), .B1(n26199), .B2(n25913), .ZN(
        n21043) );
  OAI22_X2 U1444 ( .A1(n19988), .A2(n25914), .B1(n26198), .B2(n25913), .ZN(
        n21044) );
  OAI22_X2 U1445 ( .A1(n19923), .A2(n25914), .B1(n26197), .B2(n25913), .ZN(
        n21045) );
  OAI22_X2 U1446 ( .A1(n19858), .A2(n25914), .B1(n26196), .B2(n25913), .ZN(
        n21046) );
  OAI22_X2 U1447 ( .A1(n19793), .A2(n25914), .B1(n26195), .B2(n25913), .ZN(
        n21047) );
  OAI22_X2 U1448 ( .A1(n19728), .A2(n25914), .B1(n26194), .B2(n25913), .ZN(
        n21048) );
  OAI22_X2 U1449 ( .A1(n19663), .A2(n25914), .B1(n26193), .B2(n24888), .ZN(
        n21049) );
  OAI22_X2 U1450 ( .A1(n19598), .A2(n25914), .B1(n26192), .B2(n24888), .ZN(
        n21050) );
  OAI22_X2 U1456 ( .A1(n20244), .A2(n25911), .B1(n26217), .B2(n25910), .ZN(
        n21056) );
  OAI22_X2 U1457 ( .A1(n20179), .A2(n25911), .B1(n26216), .B2(n25910), .ZN(
        n21057) );
  OAI22_X2 U1458 ( .A1(n20114), .A2(n25911), .B1(n26215), .B2(n25910), .ZN(
        n21058) );
  OAI22_X2 U1459 ( .A1(n20049), .A2(n25911), .B1(n26214), .B2(n24835), .ZN(
        n21059) );
  OAI22_X2 U1460 ( .A1(n19984), .A2(n25911), .B1(n26213), .B2(n24835), .ZN(
        n21060) );
  OAI22_X2 U1461 ( .A1(n19919), .A2(n25911), .B1(n26212), .B2(n24835), .ZN(
        n21061) );
  OAI22_X2 U1462 ( .A1(n19854), .A2(n25911), .B1(n26211), .B2(n24835), .ZN(
        n21062) );
  OAI22_X2 U1463 ( .A1(n19789), .A2(n25911), .B1(n26210), .B2(n24835), .ZN(
        n21063) );
  OAI22_X2 U1464 ( .A1(n19724), .A2(n25911), .B1(n26209), .B2(n25910), .ZN(
        n21064) );
  OAI22_X2 U1465 ( .A1(n19659), .A2(n25911), .B1(n26208), .B2(n24835), .ZN(
        n21065) );
  OAI22_X2 U1466 ( .A1(n19594), .A2(n25911), .B1(n26207), .B2(n24835), .ZN(
        n21066) );
  OAI22_X2 U1468 ( .A1(n20501), .A2(n25911), .B1(n26266), .B2(n24835), .ZN(
        n21068) );
  OAI22_X2 U1469 ( .A1(n20435), .A2(n25911), .B1(n26265), .B2(n24835), .ZN(
        n21069) );
  OAI22_X2 U1470 ( .A1(n20370), .A2(n25911), .B1(n26264), .B2(n24835), .ZN(
        n21070) );
  OAI22_X2 U1471 ( .A1(n20305), .A2(n25911), .B1(n26263), .B2(n25910), .ZN(
        n21071) );
  OAI22_X2 U1472 ( .A1(n20240), .A2(n25911), .B1(n26262), .B2(n25910), .ZN(
        n21072) );
  OAI22_X2 U1473 ( .A1(n20175), .A2(n25911), .B1(n26261), .B2(n25910), .ZN(
        n21073) );
  OAI22_X2 U1474 ( .A1(n20110), .A2(n25911), .B1(n26260), .B2(n25910), .ZN(
        n21074) );
  OAI22_X2 U1475 ( .A1(n20045), .A2(n25911), .B1(n26259), .B2(n25910), .ZN(
        n21075) );
  OAI22_X2 U1476 ( .A1(n19980), .A2(n25911), .B1(n26258), .B2(n25910), .ZN(
        n21076) );
  OAI22_X2 U1477 ( .A1(n19915), .A2(n25911), .B1(n26257), .B2(n25910), .ZN(
        n21077) );
  OAI22_X2 U1478 ( .A1(n19850), .A2(n25911), .B1(n26256), .B2(n25910), .ZN(
        n21078) );
  OAI22_X2 U1479 ( .A1(n19785), .A2(n25911), .B1(n26255), .B2(n24835), .ZN(
        n21079) );
  OAI22_X2 U1480 ( .A1(n19720), .A2(n25911), .B1(n26254), .B2(n25910), .ZN(
        n21080) );
  OAI22_X2 U1481 ( .A1(n19655), .A2(n25911), .B1(n26253), .B2(n24835), .ZN(
        n21081) );
  OAI22_X2 U1482 ( .A1(n19590), .A2(n25911), .B1(n26252), .B2(n24835), .ZN(
        n21082) );
  OAI22_X2 U1484 ( .A1(n22402), .A2(n26281), .B1(n24887), .B2(n11399), .ZN(
        n21084) );
  OAI22_X2 U1486 ( .A1(n16404), .A2(n26359), .B1(n11402), .B2(n25783), .ZN(
        n21085) );
  OAI22_X2 U1487 ( .A1(n16441), .A2(n26359), .B1(n11402), .B2(n25786), .ZN(
        n21086) );
  OAI22_X2 U1488 ( .A1(n16478), .A2(n26359), .B1(n11402), .B2(n25789), .ZN(
        n21087) );
  OAI22_X2 U1489 ( .A1(n16515), .A2(n26359), .B1(n11402), .B2(n25794), .ZN(
        n21088) );
  OAI22_X2 U1490 ( .A1(n16552), .A2(n26359), .B1(n11402), .B2(n25799), .ZN(
        n21089) );
  OAI22_X2 U1491 ( .A1(n16589), .A2(n26359), .B1(n11402), .B2(n25801), .ZN(
        n21090) );
  OAI22_X2 U1492 ( .A1(n16626), .A2(n26359), .B1(n11402), .B2(n25804), .ZN(
        n21091) );
  OAI22_X2 U1493 ( .A1(n16663), .A2(n26359), .B1(n11402), .B2(n25807), .ZN(
        n21092) );
  OAI22_X2 U1494 ( .A1(n16700), .A2(n26359), .B1(n11402), .B2(n25810), .ZN(
        n21093) );
  OAI22_X2 U1495 ( .A1(n16737), .A2(n26359), .B1(n11402), .B2(n25813), .ZN(
        n21094) );
  OAI22_X2 U1496 ( .A1(n16774), .A2(n26359), .B1(n11402), .B2(n25816), .ZN(
        n21095) );
  OAI22_X2 U1497 ( .A1(n16811), .A2(n26359), .B1(n11402), .B2(n25819), .ZN(
        n21096) );
  OAI22_X2 U1498 ( .A1(n16848), .A2(n26359), .B1(n11402), .B2(n25822), .ZN(
        n21097) );
  OAI22_X2 U1499 ( .A1(n16885), .A2(n26359), .B1(n11402), .B2(n25825), .ZN(
        n21098) );
  OAI22_X2 U1500 ( .A1(n16922), .A2(n26359), .B1(n11402), .B2(n25830), .ZN(
        n21099) );
  OAI22_X2 U1501 ( .A1(n16959), .A2(n26359), .B1(n11402), .B2(n25833), .ZN(
        n21100) );
  OAI22_X2 U1504 ( .A1(n16405), .A2(n26358), .B1(n25782), .B2(n11422), .ZN(
        n21101) );
  OAI22_X2 U1505 ( .A1(n16442), .A2(n26358), .B1(n25785), .B2(n11422), .ZN(
        n21102) );
  OAI22_X2 U1506 ( .A1(n16479), .A2(n26358), .B1(n25788), .B2(n11422), .ZN(
        n21103) );
  OAI22_X2 U1507 ( .A1(n16516), .A2(n26358), .B1(n25791), .B2(n11422), .ZN(
        n21104) );
  OAI22_X2 U1508 ( .A1(n16553), .A2(n26358), .B1(n25796), .B2(n11422), .ZN(
        n21105) );
  OAI22_X2 U1509 ( .A1(n16590), .A2(n26358), .B1(n25800), .B2(n11422), .ZN(
        n21106) );
  OAI22_X2 U1510 ( .A1(n16627), .A2(n26358), .B1(n25803), .B2(n11422), .ZN(
        n21107) );
  OAI22_X2 U1511 ( .A1(n16664), .A2(n26358), .B1(n25806), .B2(n11422), .ZN(
        n21108) );
  OAI22_X2 U1512 ( .A1(n16701), .A2(n26358), .B1(n25809), .B2(n11422), .ZN(
        n21109) );
  OAI22_X2 U1513 ( .A1(n16738), .A2(n26358), .B1(n25812), .B2(n11422), .ZN(
        n21110) );
  OAI22_X2 U1514 ( .A1(n16775), .A2(n26358), .B1(n25815), .B2(n11422), .ZN(
        n21111) );
  OAI22_X2 U1515 ( .A1(n16812), .A2(n26358), .B1(n25818), .B2(n11422), .ZN(
        n21112) );
  OAI22_X2 U1516 ( .A1(n16849), .A2(n26358), .B1(n25821), .B2(n11422), .ZN(
        n21113) );
  OAI22_X2 U1517 ( .A1(n16886), .A2(n26358), .B1(n25824), .B2(n11422), .ZN(
        n21114) );
  OAI22_X2 U1518 ( .A1(n16923), .A2(n26358), .B1(n25827), .B2(n11422), .ZN(
        n21115) );
  OAI22_X2 U1519 ( .A1(n16960), .A2(n26358), .B1(n25832), .B2(n11422), .ZN(
        n21116) );
  OAI22_X2 U1522 ( .A1(n16409), .A2(n26357), .B1(n25784), .B2(n11425), .ZN(
        n21117) );
  OAI22_X2 U1523 ( .A1(n16446), .A2(n26357), .B1(n25787), .B2(n11425), .ZN(
        n21118) );
  OAI22_X2 U1524 ( .A1(n16483), .A2(n26357), .B1(n25790), .B2(n11425), .ZN(
        n21119) );
  OAI22_X2 U1525 ( .A1(n16520), .A2(n26357), .B1(n25794), .B2(n11425), .ZN(
        n21120) );
  OAI22_X2 U1526 ( .A1(n16557), .A2(n26357), .B1(n25799), .B2(n11425), .ZN(
        n21121) );
  OAI22_X2 U1527 ( .A1(n16594), .A2(n26357), .B1(n25802), .B2(n11425), .ZN(
        n21122) );
  OAI22_X2 U1528 ( .A1(n16631), .A2(n26357), .B1(n25805), .B2(n11425), .ZN(
        n21123) );
  OAI22_X2 U1529 ( .A1(n16668), .A2(n26357), .B1(n25808), .B2(n11425), .ZN(
        n21124) );
  OAI22_X2 U1530 ( .A1(n16705), .A2(n26357), .B1(n25811), .B2(n11425), .ZN(
        n21125) );
  OAI22_X2 U1531 ( .A1(n16742), .A2(n26357), .B1(n25814), .B2(n11425), .ZN(
        n21126) );
  OAI22_X2 U1532 ( .A1(n16779), .A2(n26357), .B1(n25817), .B2(n11425), .ZN(
        n21127) );
  OAI22_X2 U1533 ( .A1(n16816), .A2(n26357), .B1(n25820), .B2(n11425), .ZN(
        n21128) );
  OAI22_X2 U1534 ( .A1(n16853), .A2(n26357), .B1(n25823), .B2(n11425), .ZN(
        n21129) );
  OAI22_X2 U1535 ( .A1(n16890), .A2(n26357), .B1(n25826), .B2(n11425), .ZN(
        n21130) );
  OAI22_X2 U1536 ( .A1(n16927), .A2(n26357), .B1(n25830), .B2(n11425), .ZN(
        n21131) );
  OAI22_X2 U1537 ( .A1(n16964), .A2(n26357), .B1(n25834), .B2(n11425), .ZN(
        n21132) );
  OAI22_X2 U1540 ( .A1(n16410), .A2(n26356), .B1(n25782), .B2(n11428), .ZN(
        n21133) );
  OAI22_X2 U1541 ( .A1(n16447), .A2(n26356), .B1(n25785), .B2(n11428), .ZN(
        n21134) );
  OAI22_X2 U1542 ( .A1(n16484), .A2(n26356), .B1(n25788), .B2(n11428), .ZN(
        n21135) );
  OAI22_X2 U1543 ( .A1(n16521), .A2(n26356), .B1(n25791), .B2(n11428), .ZN(
        n21136) );
  OAI22_X2 U1544 ( .A1(n16558), .A2(n26356), .B1(n25796), .B2(n11428), .ZN(
        n21137) );
  OAI22_X2 U1545 ( .A1(n16595), .A2(n26356), .B1(n25800), .B2(n11428), .ZN(
        n21138) );
  OAI22_X2 U1546 ( .A1(n16632), .A2(n26356), .B1(n25803), .B2(n11428), .ZN(
        n21139) );
  OAI22_X2 U1547 ( .A1(n16669), .A2(n26356), .B1(n25806), .B2(n11428), .ZN(
        n21140) );
  OAI22_X2 U1548 ( .A1(n16706), .A2(n26356), .B1(n25809), .B2(n11428), .ZN(
        n21141) );
  OAI22_X2 U1549 ( .A1(n16743), .A2(n26356), .B1(n25812), .B2(n11428), .ZN(
        n21142) );
  OAI22_X2 U1550 ( .A1(n16780), .A2(n26356), .B1(n25815), .B2(n11428), .ZN(
        n21143) );
  OAI22_X2 U1551 ( .A1(n16817), .A2(n26356), .B1(n25818), .B2(n11428), .ZN(
        n21144) );
  OAI22_X2 U1552 ( .A1(n16854), .A2(n26356), .B1(n25821), .B2(n11428), .ZN(
        n21145) );
  OAI22_X2 U1553 ( .A1(n16891), .A2(n26356), .B1(n25824), .B2(n11428), .ZN(
        n21146) );
  OAI22_X2 U1554 ( .A1(n16928), .A2(n26356), .B1(n25827), .B2(n11428), .ZN(
        n21147) );
  OAI22_X2 U1555 ( .A1(n16965), .A2(n26356), .B1(n25832), .B2(n11428), .ZN(
        n21148) );
  OAI22_X2 U1559 ( .A1(n19350), .A2(n26304), .B1(n11433), .B2(n11434), .ZN(
        n21150) );
  OAI22_X2 U1560 ( .A1(n19351), .A2(n26304), .B1(n11433), .B2(n11434), .ZN(
        n21151) );
  NAND2_X2 U1565 ( .A1(U4_DATA1_7), .A2(n25959), .ZN(n11438) );
  NAND2_X2 U1567 ( .A1(U4_DATA1_8), .A2(n25959), .ZN(n11439) );
  NAND2_X2 U1569 ( .A1(U4_DATA1_9), .A2(n25959), .ZN(n11440) );
  OAI22_X2 U1570 ( .A1(n22412), .A2(n11441), .B1(n26280), .B2(n27813), .ZN(
        n21155) );
  OAI22_X2 U1572 ( .A1(n22411), .A2(n11441), .B1(n26280), .B2(n27812), .ZN(
        n21156) );
  OAI22_X2 U1574 ( .A1(n22410), .A2(n11441), .B1(n26280), .B2(n27811), .ZN(
        n21157) );
  OAI22_X2 U1576 ( .A1(n22409), .A2(n11441), .B1(n26280), .B2(n27810), .ZN(
        n21158) );
  OAI22_X2 U1578 ( .A1(n22408), .A2(n11441), .B1(n26280), .B2(n27809), .ZN(
        n21159) );
  OAI22_X2 U1580 ( .A1(n25775), .A2(n11441), .B1(n26280), .B2(n27808), .ZN(
        n21160) );
  OAI22_X2 U1582 ( .A1(n18744), .A2(n11441), .B1(n26280), .B2(n27807), .ZN(
        n21161) );
  OAI22_X2 U1584 ( .A1(n18745), .A2(n11441), .B1(n26280), .B2(n27806), .ZN(
        n21162) );
  OAI22_X2 U1586 ( .A1(n19313), .A2(n26341), .B1(n26268), .B2(n11452), .ZN(
        n21163) );
  OAI22_X2 U1587 ( .A1(n19276), .A2(n26341), .B1(n26269), .B2(n11452), .ZN(
        n21164) );
  OAI22_X2 U1588 ( .A1(n19239), .A2(n26341), .B1(n26270), .B2(n11452), .ZN(
        n21165) );
  OAI22_X2 U1589 ( .A1(n19202), .A2(n26341), .B1(n26271), .B2(n11452), .ZN(
        n21166) );
  OAI22_X2 U1590 ( .A1(n19165), .A2(n26341), .B1(n26272), .B2(n11452), .ZN(
        n21167) );
  OAI22_X2 U1591 ( .A1(n19128), .A2(n26341), .B1(n26273), .B2(n11452), .ZN(
        n21168) );
  OAI22_X2 U1592 ( .A1(n19091), .A2(n26341), .B1(n26274), .B2(n11452), .ZN(
        n21169) );
  OAI22_X2 U1593 ( .A1(n19054), .A2(n26341), .B1(n26275), .B2(n11452), .ZN(
        n21170) );
  OAI22_X2 U1594 ( .A1(n19017), .A2(n26341), .B1(n26276), .B2(n11452), .ZN(
        n21171) );
  OAI22_X2 U1595 ( .A1(n18980), .A2(n26341), .B1(n26277), .B2(n11452), .ZN(
        n21172) );
  OAI22_X2 U1596 ( .A1(n18943), .A2(n26341), .B1(n26278), .B2(n11452), .ZN(
        n21173) );
  OAI22_X2 U1597 ( .A1(n18906), .A2(n26341), .B1(n26279), .B2(n11452), .ZN(
        n21174) );
  OAI22_X2 U1598 ( .A1(n18869), .A2(n26341), .B1(n26131), .B2(n11452), .ZN(
        n21175) );
  OAI22_X2 U1599 ( .A1(n18832), .A2(n26341), .B1(n26132), .B2(n11452), .ZN(
        n21176) );
  OAI22_X2 U1600 ( .A1(n18795), .A2(n26341), .B1(n26133), .B2(n11452), .ZN(
        n21177) );
  OAI22_X2 U1601 ( .A1(n18758), .A2(n26341), .B1(n26134), .B2(n11452), .ZN(
        n21178) );
  OAI22_X2 U1604 ( .A1(n19314), .A2(n26340), .B1(n26268), .B2(n11455), .ZN(
        n21179) );
  OAI22_X2 U1605 ( .A1(n19277), .A2(n26340), .B1(n26269), .B2(n11455), .ZN(
        n21180) );
  OAI22_X2 U1606 ( .A1(n19240), .A2(n26340), .B1(n26270), .B2(n11455), .ZN(
        n21181) );
  OAI22_X2 U1607 ( .A1(n19203), .A2(n26340), .B1(n26271), .B2(n11455), .ZN(
        n21182) );
  OAI22_X2 U1608 ( .A1(n19166), .A2(n26340), .B1(n26272), .B2(n11455), .ZN(
        n21183) );
  OAI22_X2 U1609 ( .A1(n19129), .A2(n26340), .B1(n26273), .B2(n11455), .ZN(
        n21184) );
  OAI22_X2 U1610 ( .A1(n19092), .A2(n26340), .B1(n26274), .B2(n11455), .ZN(
        n21185) );
  OAI22_X2 U1611 ( .A1(n19055), .A2(n26340), .B1(n26275), .B2(n11455), .ZN(
        n21186) );
  OAI22_X2 U1612 ( .A1(n19018), .A2(n26340), .B1(n26276), .B2(n11455), .ZN(
        n21187) );
  OAI22_X2 U1613 ( .A1(n18981), .A2(n26340), .B1(n26277), .B2(n11455), .ZN(
        n21188) );
  OAI22_X2 U1614 ( .A1(n18944), .A2(n26340), .B1(n26278), .B2(n11455), .ZN(
        n21189) );
  OAI22_X2 U1615 ( .A1(n18907), .A2(n26340), .B1(n26279), .B2(n11455), .ZN(
        n21190) );
  OAI22_X2 U1616 ( .A1(n18870), .A2(n26340), .B1(n26131), .B2(n11455), .ZN(
        n21191) );
  OAI22_X2 U1617 ( .A1(n18833), .A2(n26340), .B1(n26132), .B2(n11455), .ZN(
        n21192) );
  OAI22_X2 U1618 ( .A1(n18796), .A2(n26340), .B1(n26133), .B2(n11455), .ZN(
        n21193) );
  OAI22_X2 U1619 ( .A1(n18759), .A2(n26340), .B1(n26134), .B2(n11455), .ZN(
        n21194) );
  OAI22_X2 U1622 ( .A1(n19318), .A2(n26339), .B1(n26268), .B2(n11457), .ZN(
        n21195) );
  OAI22_X2 U1623 ( .A1(n19281), .A2(n26339), .B1(n26269), .B2(n11457), .ZN(
        n21196) );
  OAI22_X2 U1624 ( .A1(n19244), .A2(n26339), .B1(n26270), .B2(n11457), .ZN(
        n21197) );
  OAI22_X2 U1625 ( .A1(n19207), .A2(n26339), .B1(n26271), .B2(n11457), .ZN(
        n21198) );
  OAI22_X2 U1626 ( .A1(n19170), .A2(n26339), .B1(n26272), .B2(n11457), .ZN(
        n21199) );
  OAI22_X2 U1627 ( .A1(n19133), .A2(n26339), .B1(n26273), .B2(n11457), .ZN(
        n21200) );
  OAI22_X2 U1628 ( .A1(n19096), .A2(n26339), .B1(n26274), .B2(n11457), .ZN(
        n21201) );
  OAI22_X2 U1629 ( .A1(n19059), .A2(n26339), .B1(n26275), .B2(n11457), .ZN(
        n21202) );
  OAI22_X2 U1630 ( .A1(n19022), .A2(n26339), .B1(n26276), .B2(n11457), .ZN(
        n21203) );
  OAI22_X2 U1631 ( .A1(n18985), .A2(n26339), .B1(n26277), .B2(n11457), .ZN(
        n21204) );
  OAI22_X2 U1632 ( .A1(n18948), .A2(n26339), .B1(n26278), .B2(n11457), .ZN(
        n21205) );
  OAI22_X2 U1633 ( .A1(n18911), .A2(n26339), .B1(n26279), .B2(n11457), .ZN(
        n21206) );
  OAI22_X2 U1634 ( .A1(n18874), .A2(n26339), .B1(n26131), .B2(n11457), .ZN(
        n21207) );
  OAI22_X2 U1635 ( .A1(n18837), .A2(n26339), .B1(n26132), .B2(n11457), .ZN(
        n21208) );
  OAI22_X2 U1636 ( .A1(n18800), .A2(n26339), .B1(n26133), .B2(n11457), .ZN(
        n21209) );
  OAI22_X2 U1637 ( .A1(n18763), .A2(n26339), .B1(n26134), .B2(n11457), .ZN(
        n21210) );
  OAI22_X2 U1640 ( .A1(n19319), .A2(n26338), .B1(n26268), .B2(n11459), .ZN(
        n21211) );
  OAI22_X2 U1641 ( .A1(n19282), .A2(n26338), .B1(n26269), .B2(n11459), .ZN(
        n21212) );
  OAI22_X2 U1642 ( .A1(n19245), .A2(n26338), .B1(n26270), .B2(n11459), .ZN(
        n21213) );
  OAI22_X2 U1643 ( .A1(n19208), .A2(n26338), .B1(n26271), .B2(n11459), .ZN(
        n21214) );
  OAI22_X2 U1644 ( .A1(n19171), .A2(n26338), .B1(n26272), .B2(n11459), .ZN(
        n21215) );
  OAI22_X2 U1645 ( .A1(n19134), .A2(n26338), .B1(n26273), .B2(n11459), .ZN(
        n21216) );
  OAI22_X2 U1646 ( .A1(n19097), .A2(n26338), .B1(n26274), .B2(n11459), .ZN(
        n21217) );
  OAI22_X2 U1647 ( .A1(n19060), .A2(n26338), .B1(n26275), .B2(n11459), .ZN(
        n21218) );
  OAI22_X2 U1648 ( .A1(n19023), .A2(n26338), .B1(n26276), .B2(n11459), .ZN(
        n21219) );
  OAI22_X2 U1649 ( .A1(n18986), .A2(n26338), .B1(n26277), .B2(n11459), .ZN(
        n21220) );
  OAI22_X2 U1650 ( .A1(n18949), .A2(n26338), .B1(n26278), .B2(n11459), .ZN(
        n21221) );
  OAI22_X2 U1651 ( .A1(n18912), .A2(n26338), .B1(n26279), .B2(n11459), .ZN(
        n21222) );
  OAI22_X2 U1652 ( .A1(n18875), .A2(n26338), .B1(n26131), .B2(n11459), .ZN(
        n21223) );
  OAI22_X2 U1653 ( .A1(n18838), .A2(n26338), .B1(n26132), .B2(n11459), .ZN(
        n21224) );
  OAI22_X2 U1654 ( .A1(n18801), .A2(n26338), .B1(n26133), .B2(n11459), .ZN(
        n21225) );
  OAI22_X2 U1655 ( .A1(n18764), .A2(n26338), .B1(n26134), .B2(n11459), .ZN(
        n21226) );
  OAI22_X2 U1658 ( .A1(n19322), .A2(n26332), .B1(n26268), .B2(n11461), .ZN(
        n21227) );
  OAI22_X2 U1659 ( .A1(n19285), .A2(n26332), .B1(n26269), .B2(n11461), .ZN(
        n21228) );
  OAI22_X2 U1660 ( .A1(n19248), .A2(n26332), .B1(n26270), .B2(n11461), .ZN(
        n21229) );
  OAI22_X2 U1661 ( .A1(n19211), .A2(n26332), .B1(n26271), .B2(n11461), .ZN(
        n21230) );
  OAI22_X2 U1662 ( .A1(n19174), .A2(n26332), .B1(n26272), .B2(n11461), .ZN(
        n21231) );
  OAI22_X2 U1663 ( .A1(n19137), .A2(n26332), .B1(n26273), .B2(n11461), .ZN(
        n21232) );
  OAI22_X2 U1664 ( .A1(n19100), .A2(n26332), .B1(n26274), .B2(n11461), .ZN(
        n21233) );
  OAI22_X2 U1665 ( .A1(n19063), .A2(n26332), .B1(n26275), .B2(n11461), .ZN(
        n21234) );
  OAI22_X2 U1666 ( .A1(n19026), .A2(n26332), .B1(n26276), .B2(n11461), .ZN(
        n21235) );
  OAI22_X2 U1667 ( .A1(n18989), .A2(n26332), .B1(n26277), .B2(n11461), .ZN(
        n21236) );
  OAI22_X2 U1668 ( .A1(n18952), .A2(n26332), .B1(n26278), .B2(n11461), .ZN(
        n21237) );
  OAI22_X2 U1669 ( .A1(n18915), .A2(n26332), .B1(n26279), .B2(n11461), .ZN(
        n21238) );
  OAI22_X2 U1670 ( .A1(n18878), .A2(n26332), .B1(n26131), .B2(n11461), .ZN(
        n21239) );
  OAI22_X2 U1671 ( .A1(n18841), .A2(n26332), .B1(n26132), .B2(n11461), .ZN(
        n21240) );
  OAI22_X2 U1672 ( .A1(n18804), .A2(n26332), .B1(n26133), .B2(n11461), .ZN(
        n21241) );
  OAI22_X2 U1673 ( .A1(n18767), .A2(n26332), .B1(n26134), .B2(n11461), .ZN(
        n21242) );
  OAI22_X2 U1676 ( .A1(n19323), .A2(n26331), .B1(n26268), .B2(n11464), .ZN(
        n21243) );
  OAI22_X2 U1677 ( .A1(n19286), .A2(n26331), .B1(n26269), .B2(n11464), .ZN(
        n21244) );
  OAI22_X2 U1678 ( .A1(n19249), .A2(n26331), .B1(n26270), .B2(n11464), .ZN(
        n21245) );
  OAI22_X2 U1679 ( .A1(n19212), .A2(n26331), .B1(n26271), .B2(n11464), .ZN(
        n21246) );
  OAI22_X2 U1680 ( .A1(n19175), .A2(n26331), .B1(n26272), .B2(n11464), .ZN(
        n21247) );
  OAI22_X2 U1681 ( .A1(n19138), .A2(n26331), .B1(n26273), .B2(n11464), .ZN(
        n21248) );
  OAI22_X2 U1682 ( .A1(n19101), .A2(n26331), .B1(n26274), .B2(n11464), .ZN(
        n21249) );
  OAI22_X2 U1683 ( .A1(n19064), .A2(n26331), .B1(n26275), .B2(n11464), .ZN(
        n21250) );
  OAI22_X2 U1684 ( .A1(n19027), .A2(n26331), .B1(n26276), .B2(n11464), .ZN(
        n21251) );
  OAI22_X2 U1685 ( .A1(n18990), .A2(n26331), .B1(n26277), .B2(n11464), .ZN(
        n21252) );
  OAI22_X2 U1686 ( .A1(n18953), .A2(n26331), .B1(n26278), .B2(n11464), .ZN(
        n21253) );
  OAI22_X2 U1687 ( .A1(n18916), .A2(n26331), .B1(n26279), .B2(n11464), .ZN(
        n21254) );
  OAI22_X2 U1688 ( .A1(n18879), .A2(n26331), .B1(n26131), .B2(n11464), .ZN(
        n21255) );
  OAI22_X2 U1689 ( .A1(n18842), .A2(n26331), .B1(n26132), .B2(n11464), .ZN(
        n21256) );
  OAI22_X2 U1690 ( .A1(n18805), .A2(n26331), .B1(n26133), .B2(n11464), .ZN(
        n21257) );
  OAI22_X2 U1691 ( .A1(n18768), .A2(n26331), .B1(n26134), .B2(n11464), .ZN(
        n21258) );
  OAI22_X2 U1694 ( .A1(n19327), .A2(n26330), .B1(n26268), .B2(n11466), .ZN(
        n21259) );
  OAI22_X2 U1695 ( .A1(n19290), .A2(n26330), .B1(n26269), .B2(n11466), .ZN(
        n21260) );
  OAI22_X2 U1696 ( .A1(n19253), .A2(n26330), .B1(n26270), .B2(n11466), .ZN(
        n21261) );
  OAI22_X2 U1697 ( .A1(n19216), .A2(n26330), .B1(n26271), .B2(n11466), .ZN(
        n21262) );
  OAI22_X2 U1698 ( .A1(n19179), .A2(n26330), .B1(n26272), .B2(n11466), .ZN(
        n21263) );
  OAI22_X2 U1699 ( .A1(n19142), .A2(n26330), .B1(n26273), .B2(n11466), .ZN(
        n21264) );
  OAI22_X2 U1700 ( .A1(n19105), .A2(n26330), .B1(n26274), .B2(n11466), .ZN(
        n21265) );
  OAI22_X2 U1701 ( .A1(n19068), .A2(n26330), .B1(n26275), .B2(n11466), .ZN(
        n21266) );
  OAI22_X2 U1702 ( .A1(n19031), .A2(n26330), .B1(n26276), .B2(n11466), .ZN(
        n21267) );
  OAI22_X2 U1703 ( .A1(n18994), .A2(n26330), .B1(n26277), .B2(n11466), .ZN(
        n21268) );
  OAI22_X2 U1704 ( .A1(n18957), .A2(n26330), .B1(n26278), .B2(n11466), .ZN(
        n21269) );
  OAI22_X2 U1705 ( .A1(n18920), .A2(n26330), .B1(n26279), .B2(n11466), .ZN(
        n21270) );
  OAI22_X2 U1706 ( .A1(n18883), .A2(n26330), .B1(n26131), .B2(n11466), .ZN(
        n21271) );
  OAI22_X2 U1707 ( .A1(n18846), .A2(n26330), .B1(n26132), .B2(n11466), .ZN(
        n21272) );
  OAI22_X2 U1708 ( .A1(n18809), .A2(n26330), .B1(n26133), .B2(n11466), .ZN(
        n21273) );
  OAI22_X2 U1709 ( .A1(n18772), .A2(n26330), .B1(n26134), .B2(n11466), .ZN(
        n21274) );
  OAI22_X2 U1712 ( .A1(n19328), .A2(n26329), .B1(n26268), .B2(n11468), .ZN(
        n21275) );
  OAI22_X2 U1713 ( .A1(n19291), .A2(n26329), .B1(n26269), .B2(n11468), .ZN(
        n21276) );
  OAI22_X2 U1714 ( .A1(n19254), .A2(n26329), .B1(n26270), .B2(n11468), .ZN(
        n21277) );
  OAI22_X2 U1715 ( .A1(n19217), .A2(n26329), .B1(n26271), .B2(n11468), .ZN(
        n21278) );
  OAI22_X2 U1716 ( .A1(n19180), .A2(n26329), .B1(n26272), .B2(n11468), .ZN(
        n21279) );
  OAI22_X2 U1717 ( .A1(n19143), .A2(n26329), .B1(n26273), .B2(n11468), .ZN(
        n21280) );
  OAI22_X2 U1718 ( .A1(n19106), .A2(n26329), .B1(n26274), .B2(n11468), .ZN(
        n21281) );
  OAI22_X2 U1719 ( .A1(n19069), .A2(n26329), .B1(n26275), .B2(n11468), .ZN(
        n21282) );
  OAI22_X2 U1720 ( .A1(n19032), .A2(n26329), .B1(n26276), .B2(n11468), .ZN(
        n21283) );
  OAI22_X2 U1721 ( .A1(n18995), .A2(n26329), .B1(n26277), .B2(n11468), .ZN(
        n21284) );
  OAI22_X2 U1722 ( .A1(n18958), .A2(n26329), .B1(n26278), .B2(n11468), .ZN(
        n21285) );
  OAI22_X2 U1723 ( .A1(n18921), .A2(n26329), .B1(n26279), .B2(n11468), .ZN(
        n21286) );
  OAI22_X2 U1724 ( .A1(n18884), .A2(n26329), .B1(n26131), .B2(n11468), .ZN(
        n21287) );
  OAI22_X2 U1725 ( .A1(n18847), .A2(n26329), .B1(n26132), .B2(n11468), .ZN(
        n21288) );
  OAI22_X2 U1726 ( .A1(n18810), .A2(n26329), .B1(n26133), .B2(n11468), .ZN(
        n21289) );
  OAI22_X2 U1727 ( .A1(n18773), .A2(n26329), .B1(n26134), .B2(n11468), .ZN(
        n21290) );
  OAI22_X2 U1730 ( .A1(n19331), .A2(n26323), .B1(n26268), .B2(n11470), .ZN(
        n21291) );
  OAI22_X2 U1731 ( .A1(n19294), .A2(n26323), .B1(n26269), .B2(n11470), .ZN(
        n21292) );
  OAI22_X2 U1732 ( .A1(n19257), .A2(n26323), .B1(n26270), .B2(n11470), .ZN(
        n21293) );
  OAI22_X2 U1733 ( .A1(n19220), .A2(n26323), .B1(n26271), .B2(n11470), .ZN(
        n21294) );
  OAI22_X2 U1734 ( .A1(n19183), .A2(n26323), .B1(n26272), .B2(n11470), .ZN(
        n21295) );
  OAI22_X2 U1735 ( .A1(n19146), .A2(n26323), .B1(n26273), .B2(n11470), .ZN(
        n21296) );
  OAI22_X2 U1736 ( .A1(n19109), .A2(n26323), .B1(n26274), .B2(n11470), .ZN(
        n21297) );
  OAI22_X2 U1737 ( .A1(n19072), .A2(n26323), .B1(n26275), .B2(n11470), .ZN(
        n21298) );
  OAI22_X2 U1738 ( .A1(n19035), .A2(n26323), .B1(n26276), .B2(n11470), .ZN(
        n21299) );
  OAI22_X2 U1739 ( .A1(n18998), .A2(n26323), .B1(n26277), .B2(n11470), .ZN(
        n21300) );
  OAI22_X2 U1740 ( .A1(n18961), .A2(n26323), .B1(n26278), .B2(n11470), .ZN(
        n21301) );
  OAI22_X2 U1741 ( .A1(n18924), .A2(n26323), .B1(n26279), .B2(n11470), .ZN(
        n21302) );
  OAI22_X2 U1742 ( .A1(n18887), .A2(n26323), .B1(n26131), .B2(n11470), .ZN(
        n21303) );
  OAI22_X2 U1743 ( .A1(n18850), .A2(n26323), .B1(n26132), .B2(n11470), .ZN(
        n21304) );
  OAI22_X2 U1744 ( .A1(n18813), .A2(n26323), .B1(n26133), .B2(n11470), .ZN(
        n21305) );
  OAI22_X2 U1745 ( .A1(n18776), .A2(n26323), .B1(n26134), .B2(n11470), .ZN(
        n21306) );
  OAI22_X2 U1748 ( .A1(n19332), .A2(n26322), .B1(n26268), .B2(n11473), .ZN(
        n21307) );
  OAI22_X2 U1749 ( .A1(n19295), .A2(n26322), .B1(n26269), .B2(n11473), .ZN(
        n21308) );
  OAI22_X2 U1750 ( .A1(n19258), .A2(n26322), .B1(n26270), .B2(n11473), .ZN(
        n21309) );
  OAI22_X2 U1751 ( .A1(n19221), .A2(n26322), .B1(n26271), .B2(n11473), .ZN(
        n21310) );
  OAI22_X2 U1752 ( .A1(n19184), .A2(n26322), .B1(n26272), .B2(n11473), .ZN(
        n21311) );
  OAI22_X2 U1753 ( .A1(n19147), .A2(n26322), .B1(n26273), .B2(n11473), .ZN(
        n21312) );
  OAI22_X2 U1754 ( .A1(n19110), .A2(n26322), .B1(n26274), .B2(n11473), .ZN(
        n21313) );
  OAI22_X2 U1755 ( .A1(n19073), .A2(n26322), .B1(n26275), .B2(n11473), .ZN(
        n21314) );
  OAI22_X2 U1756 ( .A1(n19036), .A2(n26322), .B1(n26276), .B2(n11473), .ZN(
        n21315) );
  OAI22_X2 U1757 ( .A1(n18999), .A2(n26322), .B1(n26277), .B2(n11473), .ZN(
        n21316) );
  OAI22_X2 U1758 ( .A1(n18962), .A2(n26322), .B1(n26278), .B2(n11473), .ZN(
        n21317) );
  OAI22_X2 U1759 ( .A1(n18925), .A2(n26322), .B1(n26279), .B2(n11473), .ZN(
        n21318) );
  OAI22_X2 U1760 ( .A1(n18888), .A2(n26322), .B1(n26131), .B2(n11473), .ZN(
        n21319) );
  OAI22_X2 U1761 ( .A1(n18851), .A2(n26322), .B1(n26132), .B2(n11473), .ZN(
        n21320) );
  OAI22_X2 U1762 ( .A1(n18814), .A2(n26322), .B1(n26133), .B2(n11473), .ZN(
        n21321) );
  OAI22_X2 U1763 ( .A1(n18777), .A2(n26322), .B1(n26134), .B2(n11473), .ZN(
        n21322) );
  OAI22_X2 U1766 ( .A1(n19336), .A2(n26321), .B1(n26268), .B2(n11475), .ZN(
        n21323) );
  OAI22_X2 U1767 ( .A1(n19299), .A2(n26321), .B1(n26269), .B2(n11475), .ZN(
        n21324) );
  OAI22_X2 U1768 ( .A1(n19262), .A2(n26321), .B1(n26270), .B2(n11475), .ZN(
        n21325) );
  OAI22_X2 U1769 ( .A1(n19225), .A2(n26321), .B1(n26271), .B2(n11475), .ZN(
        n21326) );
  OAI22_X2 U1770 ( .A1(n19188), .A2(n26321), .B1(n26272), .B2(n11475), .ZN(
        n21327) );
  OAI22_X2 U1771 ( .A1(n19151), .A2(n26321), .B1(n26273), .B2(n11475), .ZN(
        n21328) );
  OAI22_X2 U1772 ( .A1(n19114), .A2(n26321), .B1(n26274), .B2(n11475), .ZN(
        n21329) );
  OAI22_X2 U1773 ( .A1(n19077), .A2(n26321), .B1(n26275), .B2(n11475), .ZN(
        n21330) );
  OAI22_X2 U1774 ( .A1(n19040), .A2(n26321), .B1(n26276), .B2(n11475), .ZN(
        n21331) );
  OAI22_X2 U1775 ( .A1(n19003), .A2(n26321), .B1(n26277), .B2(n11475), .ZN(
        n21332) );
  OAI22_X2 U1776 ( .A1(n18966), .A2(n26321), .B1(n26278), .B2(n11475), .ZN(
        n21333) );
  OAI22_X2 U1777 ( .A1(n18929), .A2(n26321), .B1(n26279), .B2(n11475), .ZN(
        n21334) );
  OAI22_X2 U1778 ( .A1(n18892), .A2(n26321), .B1(n26131), .B2(n11475), .ZN(
        n21335) );
  OAI22_X2 U1779 ( .A1(n18855), .A2(n26321), .B1(n26132), .B2(n11475), .ZN(
        n21336) );
  OAI22_X2 U1780 ( .A1(n18818), .A2(n26321), .B1(n26133), .B2(n11475), .ZN(
        n21337) );
  OAI22_X2 U1781 ( .A1(n18781), .A2(n26321), .B1(n26134), .B2(n11475), .ZN(
        n21338) );
  OAI22_X2 U1784 ( .A1(n19337), .A2(n26320), .B1(n26268), .B2(n11477), .ZN(
        n21339) );
  OAI22_X2 U1785 ( .A1(n19300), .A2(n26320), .B1(n26269), .B2(n11477), .ZN(
        n21340) );
  OAI22_X2 U1786 ( .A1(n19263), .A2(n26320), .B1(n26270), .B2(n11477), .ZN(
        n21341) );
  OAI22_X2 U1787 ( .A1(n19226), .A2(n26320), .B1(n26271), .B2(n11477), .ZN(
        n21342) );
  OAI22_X2 U1788 ( .A1(n19189), .A2(n26320), .B1(n26272), .B2(n11477), .ZN(
        n21343) );
  OAI22_X2 U1789 ( .A1(n19152), .A2(n26320), .B1(n26273), .B2(n11477), .ZN(
        n21344) );
  OAI22_X2 U1790 ( .A1(n19115), .A2(n26320), .B1(n26274), .B2(n11477), .ZN(
        n21345) );
  OAI22_X2 U1791 ( .A1(n19078), .A2(n26320), .B1(n26275), .B2(n11477), .ZN(
        n21346) );
  OAI22_X2 U1792 ( .A1(n19041), .A2(n26320), .B1(n26276), .B2(n11477), .ZN(
        n21347) );
  OAI22_X2 U1793 ( .A1(n19004), .A2(n26320), .B1(n26277), .B2(n11477), .ZN(
        n21348) );
  OAI22_X2 U1794 ( .A1(n18967), .A2(n26320), .B1(n26278), .B2(n11477), .ZN(
        n21349) );
  OAI22_X2 U1795 ( .A1(n18930), .A2(n26320), .B1(n26279), .B2(n11477), .ZN(
        n21350) );
  OAI22_X2 U1796 ( .A1(n18893), .A2(n26320), .B1(n26131), .B2(n11477), .ZN(
        n21351) );
  OAI22_X2 U1797 ( .A1(n18856), .A2(n26320), .B1(n26132), .B2(n11477), .ZN(
        n21352) );
  OAI22_X2 U1798 ( .A1(n18819), .A2(n26320), .B1(n26133), .B2(n11477), .ZN(
        n21353) );
  OAI22_X2 U1799 ( .A1(n18782), .A2(n26320), .B1(n26134), .B2(n11477), .ZN(
        n21354) );
  OAI22_X2 U1802 ( .A1(n19340), .A2(n26314), .B1(n26268), .B2(n11479), .ZN(
        n21355) );
  OAI22_X2 U1803 ( .A1(n19303), .A2(n26314), .B1(n26269), .B2(n11479), .ZN(
        n21356) );
  OAI22_X2 U1804 ( .A1(n19266), .A2(n26314), .B1(n26270), .B2(n11479), .ZN(
        n21357) );
  OAI22_X2 U1805 ( .A1(n19229), .A2(n26314), .B1(n26271), .B2(n11479), .ZN(
        n21358) );
  OAI22_X2 U1806 ( .A1(n19192), .A2(n26314), .B1(n26272), .B2(n11479), .ZN(
        n21359) );
  OAI22_X2 U1807 ( .A1(n19155), .A2(n26314), .B1(n26273), .B2(n11479), .ZN(
        n21360) );
  OAI22_X2 U1808 ( .A1(n19118), .A2(n26314), .B1(n26274), .B2(n11479), .ZN(
        n21361) );
  OAI22_X2 U1809 ( .A1(n19081), .A2(n26314), .B1(n26275), .B2(n11479), .ZN(
        n21362) );
  OAI22_X2 U1810 ( .A1(n19044), .A2(n26314), .B1(n26276), .B2(n11479), .ZN(
        n21363) );
  OAI22_X2 U1811 ( .A1(n19007), .A2(n26314), .B1(n26277), .B2(n11479), .ZN(
        n21364) );
  OAI22_X2 U1812 ( .A1(n18970), .A2(n26314), .B1(n26278), .B2(n11479), .ZN(
        n21365) );
  OAI22_X2 U1813 ( .A1(n18933), .A2(n26314), .B1(n26279), .B2(n11479), .ZN(
        n21366) );
  OAI22_X2 U1814 ( .A1(n18896), .A2(n26314), .B1(n26131), .B2(n11479), .ZN(
        n21367) );
  OAI22_X2 U1815 ( .A1(n18859), .A2(n26314), .B1(n26132), .B2(n11479), .ZN(
        n21368) );
  OAI22_X2 U1816 ( .A1(n18822), .A2(n26314), .B1(n26133), .B2(n11479), .ZN(
        n21369) );
  OAI22_X2 U1817 ( .A1(n18785), .A2(n26314), .B1(n26134), .B2(n11479), .ZN(
        n21370) );
  OAI22_X2 U1820 ( .A1(n19341), .A2(n26313), .B1(n26268), .B2(n11482), .ZN(
        n21371) );
  OAI22_X2 U1821 ( .A1(n19304), .A2(n26313), .B1(n26269), .B2(n11482), .ZN(
        n21372) );
  OAI22_X2 U1822 ( .A1(n19267), .A2(n26313), .B1(n26270), .B2(n11482), .ZN(
        n21373) );
  OAI22_X2 U1823 ( .A1(n19230), .A2(n26313), .B1(n26271), .B2(n11482), .ZN(
        n21374) );
  OAI22_X2 U1824 ( .A1(n19193), .A2(n26313), .B1(n26272), .B2(n11482), .ZN(
        n21375) );
  OAI22_X2 U1825 ( .A1(n19156), .A2(n26313), .B1(n26273), .B2(n11482), .ZN(
        n21376) );
  OAI22_X2 U1826 ( .A1(n19119), .A2(n26313), .B1(n26274), .B2(n11482), .ZN(
        n21377) );
  OAI22_X2 U1827 ( .A1(n19082), .A2(n26313), .B1(n26275), .B2(n11482), .ZN(
        n21378) );
  OAI22_X2 U1828 ( .A1(n19045), .A2(n26313), .B1(n26276), .B2(n11482), .ZN(
        n21379) );
  OAI22_X2 U1829 ( .A1(n19008), .A2(n26313), .B1(n26277), .B2(n11482), .ZN(
        n21380) );
  OAI22_X2 U1830 ( .A1(n18971), .A2(n26313), .B1(n26278), .B2(n11482), .ZN(
        n21381) );
  OAI22_X2 U1831 ( .A1(n18934), .A2(n26313), .B1(n26279), .B2(n11482), .ZN(
        n21382) );
  OAI22_X2 U1832 ( .A1(n18897), .A2(n26313), .B1(n26131), .B2(n11482), .ZN(
        n21383) );
  OAI22_X2 U1833 ( .A1(n18860), .A2(n26313), .B1(n26132), .B2(n11482), .ZN(
        n21384) );
  OAI22_X2 U1834 ( .A1(n18823), .A2(n26313), .B1(n26133), .B2(n11482), .ZN(
        n21385) );
  OAI22_X2 U1835 ( .A1(n18786), .A2(n26313), .B1(n26134), .B2(n11482), .ZN(
        n21386) );
  OAI22_X2 U1838 ( .A1(n19345), .A2(n26312), .B1(n26268), .B2(n11484), .ZN(
        n21387) );
  OAI22_X2 U1839 ( .A1(n19308), .A2(n26312), .B1(n26269), .B2(n11484), .ZN(
        n21388) );
  OAI22_X2 U1840 ( .A1(n19271), .A2(n26312), .B1(n26270), .B2(n11484), .ZN(
        n21389) );
  OAI22_X2 U1841 ( .A1(n19234), .A2(n26312), .B1(n26271), .B2(n11484), .ZN(
        n21390) );
  OAI22_X2 U1842 ( .A1(n19197), .A2(n26312), .B1(n26272), .B2(n11484), .ZN(
        n21391) );
  OAI22_X2 U1843 ( .A1(n19160), .A2(n26312), .B1(n26273), .B2(n11484), .ZN(
        n21392) );
  OAI22_X2 U1844 ( .A1(n19123), .A2(n26312), .B1(n26274), .B2(n11484), .ZN(
        n21393) );
  OAI22_X2 U1845 ( .A1(n19086), .A2(n26312), .B1(n26275), .B2(n11484), .ZN(
        n21394) );
  OAI22_X2 U1846 ( .A1(n19049), .A2(n26312), .B1(n26276), .B2(n11484), .ZN(
        n21395) );
  OAI22_X2 U1847 ( .A1(n19012), .A2(n26312), .B1(n26277), .B2(n11484), .ZN(
        n21396) );
  OAI22_X2 U1848 ( .A1(n18975), .A2(n26312), .B1(n26278), .B2(n11484), .ZN(
        n21397) );
  OAI22_X2 U1849 ( .A1(n18938), .A2(n26312), .B1(n26279), .B2(n11484), .ZN(
        n21398) );
  OAI22_X2 U1850 ( .A1(n18901), .A2(n26312), .B1(n26131), .B2(n11484), .ZN(
        n21399) );
  OAI22_X2 U1851 ( .A1(n18864), .A2(n26312), .B1(n26132), .B2(n11484), .ZN(
        n21400) );
  OAI22_X2 U1852 ( .A1(n18827), .A2(n26312), .B1(n26133), .B2(n11484), .ZN(
        n21401) );
  OAI22_X2 U1853 ( .A1(n18790), .A2(n26312), .B1(n26134), .B2(n11484), .ZN(
        n21402) );
  OAI22_X2 U1856 ( .A1(n19346), .A2(n26311), .B1(n26268), .B2(n11486), .ZN(
        n21403) );
  OAI22_X2 U1857 ( .A1(n19309), .A2(n26311), .B1(n26269), .B2(n11486), .ZN(
        n21404) );
  OAI22_X2 U1858 ( .A1(n19272), .A2(n26311), .B1(n26270), .B2(n11486), .ZN(
        n21405) );
  OAI22_X2 U1859 ( .A1(n19235), .A2(n26311), .B1(n26271), .B2(n11486), .ZN(
        n21406) );
  OAI22_X2 U1860 ( .A1(n19198), .A2(n26311), .B1(n26272), .B2(n11486), .ZN(
        n21407) );
  OAI22_X2 U1861 ( .A1(n19161), .A2(n26311), .B1(n26273), .B2(n11486), .ZN(
        n21408) );
  OAI22_X2 U1862 ( .A1(n19124), .A2(n26311), .B1(n26274), .B2(n11486), .ZN(
        n21409) );
  OAI22_X2 U1863 ( .A1(n19087), .A2(n26311), .B1(n26275), .B2(n11486), .ZN(
        n21410) );
  OAI22_X2 U1864 ( .A1(n19050), .A2(n26311), .B1(n26276), .B2(n11486), .ZN(
        n21411) );
  OAI22_X2 U1865 ( .A1(n19013), .A2(n26311), .B1(n26277), .B2(n11486), .ZN(
        n21412) );
  OAI22_X2 U1866 ( .A1(n18976), .A2(n26311), .B1(n26278), .B2(n11486), .ZN(
        n21413) );
  OAI22_X2 U1867 ( .A1(n18939), .A2(n26311), .B1(n26279), .B2(n11486), .ZN(
        n21414) );
  OAI22_X2 U1868 ( .A1(n18902), .A2(n26311), .B1(n26131), .B2(n11486), .ZN(
        n21415) );
  OAI22_X2 U1869 ( .A1(n18865), .A2(n26311), .B1(n26132), .B2(n11486), .ZN(
        n21416) );
  OAI22_X2 U1870 ( .A1(n18828), .A2(n26311), .B1(n26133), .B2(n11486), .ZN(
        n21417) );
  OAI22_X2 U1871 ( .A1(n18791), .A2(n26311), .B1(n26134), .B2(n11486), .ZN(
        n21418) );
  NAND4_X2 U1875 ( .A1(n11487), .A2(n11490), .A3(n11491), .A4(n11492), .ZN(
        n11488) );
  OAI221_X2 U1876 ( .B1(n26459), .B2(n11494), .C1(n16371), .C2(n11487), .A(
        n26461), .ZN(n21420) );
  NAND2_X2 U1878 ( .A1(n11497), .A2(n11498), .ZN(n11494) );
  OAI22_X2 U1879 ( .A1(n16395), .A2(n26470), .B1(n25783), .B2(n11500), .ZN(
        n21421) );
  OAI22_X2 U1880 ( .A1(n16432), .A2(n26470), .B1(n25786), .B2(n11500), .ZN(
        n21422) );
  OAI22_X2 U1881 ( .A1(n16469), .A2(n26470), .B1(n25789), .B2(n11500), .ZN(
        n21423) );
  OAI22_X2 U1882 ( .A1(n16506), .A2(n26470), .B1(n25792), .B2(n11500), .ZN(
        n21424) );
  OAI22_X2 U1883 ( .A1(n16543), .A2(n26470), .B1(n25797), .B2(n11500), .ZN(
        n21425) );
  OAI22_X2 U1884 ( .A1(n16580), .A2(n26470), .B1(n25801), .B2(n11500), .ZN(
        n21426) );
  OAI22_X2 U1885 ( .A1(n16617), .A2(n26470), .B1(n25804), .B2(n11500), .ZN(
        n21427) );
  OAI22_X2 U1886 ( .A1(n16654), .A2(n26470), .B1(n25807), .B2(n11500), .ZN(
        n21428) );
  OAI22_X2 U1887 ( .A1(n16691), .A2(n26470), .B1(n25810), .B2(n11500), .ZN(
        n21429) );
  OAI22_X2 U1888 ( .A1(n16728), .A2(n26470), .B1(n25813), .B2(n11500), .ZN(
        n21430) );
  OAI22_X2 U1889 ( .A1(n16765), .A2(n26470), .B1(n25816), .B2(n11500), .ZN(
        n21431) );
  OAI22_X2 U1890 ( .A1(n16802), .A2(n26470), .B1(n25819), .B2(n11500), .ZN(
        n21432) );
  OAI22_X2 U1891 ( .A1(n16839), .A2(n26470), .B1(n25822), .B2(n11500), .ZN(
        n21433) );
  OAI22_X2 U1892 ( .A1(n16876), .A2(n26470), .B1(n25825), .B2(n11500), .ZN(
        n21434) );
  OAI22_X2 U1893 ( .A1(n16913), .A2(n26470), .B1(n25828), .B2(n11500), .ZN(
        n21435) );
  OAI22_X2 U1894 ( .A1(n16950), .A2(n26470), .B1(n25833), .B2(n11500), .ZN(
        n21436) );
  OAI22_X2 U1897 ( .A1(n16396), .A2(n26469), .B1(n25784), .B2(n11503), .ZN(
        n21437) );
  OAI22_X2 U1898 ( .A1(n16433), .A2(n26469), .B1(n25787), .B2(n11503), .ZN(
        n21438) );
  OAI22_X2 U1899 ( .A1(n16470), .A2(n26469), .B1(n25790), .B2(n11503), .ZN(
        n21439) );
  OAI22_X2 U1900 ( .A1(n16507), .A2(n26469), .B1(n25795), .B2(n11503), .ZN(
        n21440) );
  OAI22_X2 U1901 ( .A1(n16544), .A2(n26469), .B1(n25797), .B2(n11503), .ZN(
        n21441) );
  OAI22_X2 U1902 ( .A1(n16581), .A2(n26469), .B1(n25802), .B2(n11503), .ZN(
        n21442) );
  OAI22_X2 U1903 ( .A1(n16618), .A2(n26469), .B1(n25805), .B2(n11503), .ZN(
        n21443) );
  OAI22_X2 U1904 ( .A1(n16655), .A2(n26469), .B1(n25808), .B2(n11503), .ZN(
        n21444) );
  OAI22_X2 U1905 ( .A1(n16692), .A2(n26469), .B1(n25811), .B2(n11503), .ZN(
        n21445) );
  OAI22_X2 U1906 ( .A1(n16729), .A2(n26469), .B1(n25814), .B2(n11503), .ZN(
        n21446) );
  OAI22_X2 U1907 ( .A1(n16766), .A2(n26469), .B1(n25817), .B2(n11503), .ZN(
        n21447) );
  OAI22_X2 U1908 ( .A1(n16803), .A2(n26469), .B1(n25820), .B2(n11503), .ZN(
        n21448) );
  OAI22_X2 U1909 ( .A1(n16840), .A2(n26469), .B1(n25823), .B2(n11503), .ZN(
        n21449) );
  OAI22_X2 U1910 ( .A1(n16877), .A2(n26469), .B1(n25826), .B2(n11503), .ZN(
        n21450) );
  OAI22_X2 U1911 ( .A1(n16914), .A2(n26469), .B1(n25831), .B2(n11503), .ZN(
        n21451) );
  OAI22_X2 U1912 ( .A1(n16951), .A2(n26469), .B1(n25834), .B2(n11503), .ZN(
        n21452) );
  OAI22_X2 U1915 ( .A1(n16400), .A2(n26468), .B1(n25782), .B2(n11505), .ZN(
        n21453) );
  OAI22_X2 U1916 ( .A1(n16437), .A2(n26468), .B1(n25785), .B2(n11505), .ZN(
        n21454) );
  OAI22_X2 U1917 ( .A1(n16474), .A2(n26468), .B1(n25788), .B2(n11505), .ZN(
        n21455) );
  OAI22_X2 U1918 ( .A1(n16511), .A2(n26468), .B1(n25794), .B2(n11505), .ZN(
        n21456) );
  OAI22_X2 U1919 ( .A1(n16548), .A2(n26468), .B1(n25799), .B2(n11505), .ZN(
        n21457) );
  OAI22_X2 U1920 ( .A1(n16585), .A2(n26468), .B1(n25800), .B2(n11505), .ZN(
        n21458) );
  OAI22_X2 U1921 ( .A1(n16622), .A2(n26468), .B1(n25803), .B2(n11505), .ZN(
        n21459) );
  OAI22_X2 U1922 ( .A1(n16659), .A2(n26468), .B1(n25806), .B2(n11505), .ZN(
        n21460) );
  OAI22_X2 U1923 ( .A1(n16696), .A2(n26468), .B1(n25809), .B2(n11505), .ZN(
        n21461) );
  OAI22_X2 U1924 ( .A1(n16733), .A2(n26468), .B1(n25812), .B2(n11505), .ZN(
        n21462) );
  OAI22_X2 U1925 ( .A1(n16770), .A2(n26468), .B1(n25815), .B2(n11505), .ZN(
        n21463) );
  OAI22_X2 U1926 ( .A1(n16807), .A2(n26468), .B1(n25818), .B2(n11505), .ZN(
        n21464) );
  OAI22_X2 U1927 ( .A1(n16844), .A2(n26468), .B1(n25821), .B2(n11505), .ZN(
        n21465) );
  OAI22_X2 U1928 ( .A1(n16881), .A2(n26468), .B1(n25824), .B2(n11505), .ZN(
        n21466) );
  OAI22_X2 U1929 ( .A1(n16918), .A2(n26468), .B1(n25830), .B2(n11505), .ZN(
        n21467) );
  OAI22_X2 U1930 ( .A1(n16955), .A2(n26468), .B1(n25832), .B2(n11505), .ZN(
        n21468) );
  OAI22_X2 U1933 ( .A1(n16401), .A2(n26467), .B1(n25783), .B2(n11507), .ZN(
        n21469) );
  OAI22_X2 U1934 ( .A1(n16438), .A2(n26467), .B1(n25786), .B2(n11507), .ZN(
        n21470) );
  OAI22_X2 U1935 ( .A1(n16475), .A2(n26467), .B1(n25789), .B2(n11507), .ZN(
        n21471) );
  OAI22_X2 U1936 ( .A1(n16512), .A2(n26467), .B1(n25795), .B2(n11507), .ZN(
        n21472) );
  OAI22_X2 U1937 ( .A1(n16549), .A2(n26467), .B1(n25796), .B2(n11507), .ZN(
        n21473) );
  OAI22_X2 U1938 ( .A1(n16586), .A2(n26467), .B1(n25801), .B2(n11507), .ZN(
        n21474) );
  OAI22_X2 U1939 ( .A1(n16623), .A2(n26467), .B1(n25804), .B2(n11507), .ZN(
        n21475) );
  OAI22_X2 U1940 ( .A1(n16660), .A2(n26467), .B1(n25807), .B2(n11507), .ZN(
        n21476) );
  OAI22_X2 U1941 ( .A1(n16697), .A2(n26467), .B1(n25810), .B2(n11507), .ZN(
        n21477) );
  OAI22_X2 U1942 ( .A1(n16734), .A2(n26467), .B1(n25813), .B2(n11507), .ZN(
        n21478) );
  OAI22_X2 U1943 ( .A1(n16771), .A2(n26467), .B1(n25816), .B2(n11507), .ZN(
        n21479) );
  OAI22_X2 U1944 ( .A1(n16808), .A2(n26467), .B1(n25819), .B2(n11507), .ZN(
        n21480) );
  OAI22_X2 U1945 ( .A1(n16845), .A2(n26467), .B1(n25822), .B2(n11507), .ZN(
        n21481) );
  OAI22_X2 U1946 ( .A1(n16882), .A2(n26467), .B1(n25825), .B2(n11507), .ZN(
        n21482) );
  OAI22_X2 U1947 ( .A1(n16919), .A2(n26467), .B1(n25831), .B2(n11507), .ZN(
        n21483) );
  OAI22_X2 U1948 ( .A1(n16956), .A2(n26467), .B1(n25833), .B2(n11507), .ZN(
        n21484) );
  OAI22_X2 U1951 ( .A1(n18171), .A2(n26479), .B1(n25784), .B2(n11509), .ZN(
        n21485) );
  OAI22_X2 U1952 ( .A1(n18208), .A2(n26479), .B1(n25787), .B2(n11509), .ZN(
        n21486) );
  OAI22_X2 U1953 ( .A1(n18245), .A2(n26479), .B1(n25790), .B2(n11509), .ZN(
        n21487) );
  OAI22_X2 U1954 ( .A1(n18282), .A2(n26479), .B1(n25791), .B2(n11509), .ZN(
        n21488) );
  OAI22_X2 U1955 ( .A1(n18319), .A2(n26479), .B1(n25796), .B2(n11509), .ZN(
        n21489) );
  OAI22_X2 U1956 ( .A1(n18356), .A2(n26479), .B1(n25802), .B2(n11509), .ZN(
        n21490) );
  OAI22_X2 U1957 ( .A1(n18393), .A2(n26479), .B1(n25805), .B2(n11509), .ZN(
        n21491) );
  OAI22_X2 U1958 ( .A1(n18430), .A2(n26479), .B1(n25808), .B2(n11509), .ZN(
        n21492) );
  OAI22_X2 U1959 ( .A1(n18467), .A2(n26479), .B1(n25811), .B2(n11509), .ZN(
        n21493) );
  OAI22_X2 U1960 ( .A1(n18504), .A2(n26479), .B1(n25814), .B2(n11509), .ZN(
        n21494) );
  OAI22_X2 U1961 ( .A1(n18541), .A2(n26479), .B1(n25817), .B2(n11509), .ZN(
        n21495) );
  OAI22_X2 U1962 ( .A1(n18578), .A2(n26479), .B1(n25820), .B2(n11509), .ZN(
        n21496) );
  OAI22_X2 U1963 ( .A1(n18615), .A2(n26479), .B1(n25823), .B2(n11509), .ZN(
        n21497) );
  OAI22_X2 U1964 ( .A1(n18652), .A2(n26479), .B1(n25826), .B2(n11509), .ZN(
        n21498) );
  OAI22_X2 U1965 ( .A1(n18689), .A2(n26479), .B1(n25827), .B2(n11509), .ZN(
        n21499) );
  OAI22_X2 U1966 ( .A1(n18726), .A2(n26479), .B1(n25834), .B2(n11509), .ZN(
        n21500) );
  OAI22_X2 U1969 ( .A1(n18172), .A2(n26478), .B1(n25782), .B2(n11512), .ZN(
        n21501) );
  OAI22_X2 U1970 ( .A1(n18209), .A2(n26478), .B1(n25785), .B2(n11512), .ZN(
        n21502) );
  OAI22_X2 U1971 ( .A1(n18246), .A2(n26478), .B1(n25788), .B2(n11512), .ZN(
        n21503) );
  OAI22_X2 U1972 ( .A1(n18283), .A2(n26478), .B1(n25792), .B2(n11512), .ZN(
        n21504) );
  OAI22_X2 U1973 ( .A1(n18320), .A2(n26478), .B1(n25797), .B2(n11512), .ZN(
        n21505) );
  OAI22_X2 U1974 ( .A1(n18357), .A2(n26478), .B1(n25800), .B2(n11512), .ZN(
        n21506) );
  OAI22_X2 U1975 ( .A1(n18394), .A2(n26478), .B1(n25803), .B2(n11512), .ZN(
        n21507) );
  OAI22_X2 U1976 ( .A1(n18431), .A2(n26478), .B1(n25806), .B2(n11512), .ZN(
        n21508) );
  OAI22_X2 U1977 ( .A1(n18468), .A2(n26478), .B1(n25809), .B2(n11512), .ZN(
        n21509) );
  OAI22_X2 U1978 ( .A1(n18505), .A2(n26478), .B1(n25812), .B2(n11512), .ZN(
        n21510) );
  OAI22_X2 U1979 ( .A1(n18542), .A2(n26478), .B1(n25815), .B2(n11512), .ZN(
        n21511) );
  OAI22_X2 U1980 ( .A1(n18579), .A2(n26478), .B1(n25818), .B2(n11512), .ZN(
        n21512) );
  OAI22_X2 U1981 ( .A1(n18616), .A2(n26478), .B1(n25821), .B2(n11512), .ZN(
        n21513) );
  OAI22_X2 U1982 ( .A1(n18653), .A2(n26478), .B1(n25824), .B2(n11512), .ZN(
        n21514) );
  OAI22_X2 U1983 ( .A1(n18690), .A2(n26478), .B1(n25828), .B2(n11512), .ZN(
        n21515) );
  OAI22_X2 U1984 ( .A1(n18727), .A2(n26478), .B1(n25832), .B2(n11512), .ZN(
        n21516) );
  OAI22_X2 U1987 ( .A1(n18176), .A2(n26477), .B1(n25784), .B2(n11514), .ZN(
        n21517) );
  OAI22_X2 U1988 ( .A1(n18213), .A2(n26477), .B1(n25787), .B2(n11514), .ZN(
        n21518) );
  OAI22_X2 U1989 ( .A1(n18250), .A2(n26477), .B1(n25790), .B2(n11514), .ZN(
        n21519) );
  OAI22_X2 U1990 ( .A1(n18287), .A2(n26477), .B1(n25795), .B2(n11514), .ZN(
        n21520) );
  OAI22_X2 U1991 ( .A1(n18324), .A2(n26477), .B1(n25799), .B2(n11514), .ZN(
        n21521) );
  OAI22_X2 U1992 ( .A1(n18361), .A2(n26477), .B1(n25802), .B2(n11514), .ZN(
        n21522) );
  OAI22_X2 U1993 ( .A1(n18398), .A2(n26477), .B1(n25805), .B2(n11514), .ZN(
        n21523) );
  OAI22_X2 U1994 ( .A1(n18435), .A2(n26477), .B1(n25808), .B2(n11514), .ZN(
        n21524) );
  OAI22_X2 U1995 ( .A1(n18472), .A2(n26477), .B1(n25811), .B2(n11514), .ZN(
        n21525) );
  OAI22_X2 U1996 ( .A1(n18509), .A2(n26477), .B1(n25814), .B2(n11514), .ZN(
        n21526) );
  OAI22_X2 U1997 ( .A1(n18546), .A2(n26477), .B1(n25817), .B2(n11514), .ZN(
        n21527) );
  OAI22_X2 U1998 ( .A1(n18583), .A2(n26477), .B1(n25820), .B2(n11514), .ZN(
        n21528) );
  OAI22_X2 U1999 ( .A1(n18620), .A2(n26477), .B1(n25823), .B2(n11514), .ZN(
        n21529) );
  OAI22_X2 U2000 ( .A1(n18657), .A2(n26477), .B1(n25826), .B2(n11514), .ZN(
        n21530) );
  OAI22_X2 U2001 ( .A1(n18694), .A2(n26477), .B1(n25831), .B2(n11514), .ZN(
        n21531) );
  OAI22_X2 U2002 ( .A1(n18731), .A2(n26477), .B1(n25834), .B2(n11514), .ZN(
        n21532) );
  OAI22_X2 U2005 ( .A1(n18177), .A2(n26476), .B1(n25783), .B2(n11516), .ZN(
        n21533) );
  OAI22_X2 U2006 ( .A1(n18214), .A2(n26476), .B1(n25786), .B2(n11516), .ZN(
        n21534) );
  OAI22_X2 U2007 ( .A1(n18251), .A2(n26476), .B1(n25789), .B2(n11516), .ZN(
        n21535) );
  OAI22_X2 U2008 ( .A1(n18288), .A2(n26476), .B1(n25794), .B2(n11516), .ZN(
        n21536) );
  OAI22_X2 U2009 ( .A1(n18325), .A2(n26476), .B1(n25799), .B2(n11516), .ZN(
        n21537) );
  OAI22_X2 U2010 ( .A1(n18362), .A2(n26476), .B1(n25801), .B2(n11516), .ZN(
        n21538) );
  OAI22_X2 U2011 ( .A1(n18399), .A2(n26476), .B1(n25804), .B2(n11516), .ZN(
        n21539) );
  OAI22_X2 U2012 ( .A1(n18436), .A2(n26476), .B1(n25807), .B2(n11516), .ZN(
        n21540) );
  OAI22_X2 U2013 ( .A1(n18473), .A2(n26476), .B1(n25810), .B2(n11516), .ZN(
        n21541) );
  OAI22_X2 U2014 ( .A1(n18510), .A2(n26476), .B1(n25813), .B2(n11516), .ZN(
        n21542) );
  OAI22_X2 U2015 ( .A1(n18547), .A2(n26476), .B1(n25816), .B2(n11516), .ZN(
        n21543) );
  OAI22_X2 U2016 ( .A1(n18584), .A2(n26476), .B1(n25819), .B2(n11516), .ZN(
        n21544) );
  OAI22_X2 U2017 ( .A1(n18621), .A2(n26476), .B1(n25822), .B2(n11516), .ZN(
        n21545) );
  OAI22_X2 U2018 ( .A1(n18658), .A2(n26476), .B1(n25825), .B2(n11516), .ZN(
        n21546) );
  OAI22_X2 U2019 ( .A1(n18695), .A2(n26476), .B1(n25830), .B2(n11516), .ZN(
        n21547) );
  OAI22_X2 U2020 ( .A1(n18732), .A2(n26476), .B1(n25833), .B2(n11516), .ZN(
        n21548) );
  OAI22_X2 U2023 ( .A1(n17579), .A2(n26488), .B1(n25782), .B2(n11518), .ZN(
        n21549) );
  OAI22_X2 U2024 ( .A1(n17616), .A2(n26488), .B1(n25785), .B2(n11518), .ZN(
        n21550) );
  OAI22_X2 U2025 ( .A1(n17653), .A2(n26488), .B1(n25788), .B2(n11518), .ZN(
        n21551) );
  OAI22_X2 U2026 ( .A1(n17690), .A2(n26488), .B1(n25791), .B2(n11518), .ZN(
        n21552) );
  OAI22_X2 U2027 ( .A1(n17727), .A2(n26488), .B1(n25796), .B2(n11518), .ZN(
        n21553) );
  OAI22_X2 U2028 ( .A1(n17764), .A2(n26488), .B1(n25800), .B2(n11518), .ZN(
        n21554) );
  OAI22_X2 U2029 ( .A1(n17801), .A2(n26488), .B1(n25803), .B2(n11518), .ZN(
        n21555) );
  OAI22_X2 U2030 ( .A1(n17838), .A2(n26488), .B1(n25806), .B2(n11518), .ZN(
        n21556) );
  OAI22_X2 U2031 ( .A1(n17875), .A2(n26488), .B1(n25809), .B2(n11518), .ZN(
        n21557) );
  OAI22_X2 U2032 ( .A1(n17912), .A2(n26488), .B1(n25812), .B2(n11518), .ZN(
        n21558) );
  OAI22_X2 U2033 ( .A1(n17949), .A2(n26488), .B1(n25815), .B2(n11518), .ZN(
        n21559) );
  OAI22_X2 U2034 ( .A1(n17986), .A2(n26488), .B1(n25818), .B2(n11518), .ZN(
        n21560) );
  OAI22_X2 U2035 ( .A1(n18023), .A2(n26488), .B1(n25821), .B2(n11518), .ZN(
        n21561) );
  OAI22_X2 U2036 ( .A1(n18060), .A2(n26488), .B1(n25824), .B2(n11518), .ZN(
        n21562) );
  OAI22_X2 U2037 ( .A1(n18097), .A2(n26488), .B1(n25827), .B2(n11518), .ZN(
        n21563) );
  OAI22_X2 U2038 ( .A1(n18134), .A2(n26488), .B1(n25832), .B2(n11518), .ZN(
        n21564) );
  OAI22_X2 U2041 ( .A1(n17580), .A2(n26487), .B1(n25784), .B2(n11521), .ZN(
        n21565) );
  OAI22_X2 U2042 ( .A1(n17617), .A2(n26487), .B1(n25787), .B2(n11521), .ZN(
        n21566) );
  OAI22_X2 U2043 ( .A1(n17654), .A2(n26487), .B1(n25790), .B2(n11521), .ZN(
        n21567) );
  OAI22_X2 U2044 ( .A1(n17691), .A2(n26487), .B1(n25791), .B2(n11521), .ZN(
        n21568) );
  OAI22_X2 U2045 ( .A1(n17728), .A2(n26487), .B1(n25796), .B2(n11521), .ZN(
        n21569) );
  OAI22_X2 U2046 ( .A1(n17765), .A2(n26487), .B1(n25802), .B2(n11521), .ZN(
        n21570) );
  OAI22_X2 U2047 ( .A1(n17802), .A2(n26487), .B1(n25805), .B2(n11521), .ZN(
        n21571) );
  OAI22_X2 U2048 ( .A1(n17839), .A2(n26487), .B1(n25808), .B2(n11521), .ZN(
        n21572) );
  OAI22_X2 U2049 ( .A1(n17876), .A2(n26487), .B1(n25811), .B2(n11521), .ZN(
        n21573) );
  OAI22_X2 U2050 ( .A1(n17913), .A2(n26487), .B1(n25814), .B2(n11521), .ZN(
        n21574) );
  OAI22_X2 U2051 ( .A1(n17950), .A2(n26487), .B1(n25817), .B2(n11521), .ZN(
        n21575) );
  OAI22_X2 U2052 ( .A1(n17987), .A2(n26487), .B1(n25820), .B2(n11521), .ZN(
        n21576) );
  OAI22_X2 U2053 ( .A1(n18024), .A2(n26487), .B1(n25823), .B2(n11521), .ZN(
        n21577) );
  OAI22_X2 U2054 ( .A1(n18061), .A2(n26487), .B1(n25826), .B2(n11521), .ZN(
        n21578) );
  OAI22_X2 U2055 ( .A1(n18098), .A2(n26487), .B1(n25827), .B2(n11521), .ZN(
        n21579) );
  OAI22_X2 U2056 ( .A1(n18135), .A2(n26487), .B1(n25834), .B2(n11521), .ZN(
        n21580) );
  OAI22_X2 U2059 ( .A1(n17584), .A2(n26486), .B1(n25783), .B2(n11523), .ZN(
        n21581) );
  OAI22_X2 U2060 ( .A1(n17621), .A2(n26486), .B1(n25786), .B2(n11523), .ZN(
        n21582) );
  OAI22_X2 U2061 ( .A1(n17658), .A2(n26486), .B1(n25789), .B2(n11523), .ZN(
        n21583) );
  OAI22_X2 U2062 ( .A1(n17695), .A2(n26486), .B1(n25791), .B2(n11523), .ZN(
        n21584) );
  OAI22_X2 U2063 ( .A1(n17732), .A2(n26486), .B1(n25796), .B2(n11523), .ZN(
        n21585) );
  OAI22_X2 U2064 ( .A1(n17769), .A2(n26486), .B1(n25801), .B2(n11523), .ZN(
        n21586) );
  OAI22_X2 U2065 ( .A1(n17806), .A2(n26486), .B1(n25804), .B2(n11523), .ZN(
        n21587) );
  OAI22_X2 U2066 ( .A1(n17843), .A2(n26486), .B1(n25807), .B2(n11523), .ZN(
        n21588) );
  OAI22_X2 U2067 ( .A1(n17880), .A2(n26486), .B1(n25810), .B2(n11523), .ZN(
        n21589) );
  OAI22_X2 U2068 ( .A1(n17917), .A2(n26486), .B1(n25813), .B2(n11523), .ZN(
        n21590) );
  OAI22_X2 U2069 ( .A1(n17954), .A2(n26486), .B1(n25816), .B2(n11523), .ZN(
        n21591) );
  OAI22_X2 U2070 ( .A1(n17991), .A2(n26486), .B1(n25819), .B2(n11523), .ZN(
        n21592) );
  OAI22_X2 U2071 ( .A1(n18028), .A2(n26486), .B1(n25822), .B2(n11523), .ZN(
        n21593) );
  OAI22_X2 U2072 ( .A1(n18065), .A2(n26486), .B1(n25825), .B2(n11523), .ZN(
        n21594) );
  OAI22_X2 U2073 ( .A1(n18102), .A2(n26486), .B1(n25827), .B2(n11523), .ZN(
        n21595) );
  OAI22_X2 U2074 ( .A1(n18139), .A2(n26486), .B1(n25833), .B2(n11523), .ZN(
        n21596) );
  OAI22_X2 U2077 ( .A1(n17585), .A2(n26485), .B1(n25783), .B2(n11525), .ZN(
        n21597) );
  OAI22_X2 U2078 ( .A1(n17622), .A2(n26485), .B1(n25786), .B2(n11525), .ZN(
        n21598) );
  OAI22_X2 U2079 ( .A1(n17659), .A2(n26485), .B1(n25789), .B2(n11525), .ZN(
        n21599) );
  OAI22_X2 U2080 ( .A1(n17696), .A2(n26485), .B1(n25792), .B2(n11525), .ZN(
        n21600) );
  OAI22_X2 U2081 ( .A1(n17733), .A2(n26485), .B1(n25797), .B2(n11525), .ZN(
        n21601) );
  OAI22_X2 U2082 ( .A1(n17770), .A2(n26485), .B1(n25801), .B2(n11525), .ZN(
        n21602) );
  OAI22_X2 U2083 ( .A1(n17807), .A2(n26485), .B1(n25804), .B2(n11525), .ZN(
        n21603) );
  OAI22_X2 U2084 ( .A1(n17844), .A2(n26485), .B1(n25807), .B2(n11525), .ZN(
        n21604) );
  OAI22_X2 U2085 ( .A1(n17881), .A2(n26485), .B1(n25810), .B2(n11525), .ZN(
        n21605) );
  OAI22_X2 U2086 ( .A1(n17918), .A2(n26485), .B1(n25813), .B2(n11525), .ZN(
        n21606) );
  OAI22_X2 U2087 ( .A1(n17955), .A2(n26485), .B1(n25816), .B2(n11525), .ZN(
        n21607) );
  OAI22_X2 U2088 ( .A1(n17992), .A2(n26485), .B1(n25819), .B2(n11525), .ZN(
        n21608) );
  OAI22_X2 U2089 ( .A1(n18029), .A2(n26485), .B1(n25822), .B2(n11525), .ZN(
        n21609) );
  OAI22_X2 U2090 ( .A1(n18066), .A2(n26485), .B1(n25825), .B2(n11525), .ZN(
        n21610) );
  OAI22_X2 U2091 ( .A1(n18103), .A2(n26485), .B1(n25828), .B2(n11525), .ZN(
        n21611) );
  OAI22_X2 U2092 ( .A1(n18140), .A2(n26485), .B1(n25833), .B2(n11525), .ZN(
        n21612) );
  OAI22_X2 U2095 ( .A1(n16987), .A2(n26497), .B1(n25782), .B2(n11527), .ZN(
        n21613) );
  OAI22_X2 U2096 ( .A1(n17024), .A2(n26497), .B1(n25785), .B2(n11527), .ZN(
        n21614) );
  OAI22_X2 U2097 ( .A1(n17061), .A2(n26497), .B1(n25788), .B2(n11527), .ZN(
        n21615) );
  OAI22_X2 U2098 ( .A1(n17098), .A2(n26497), .B1(n25795), .B2(n11527), .ZN(
        n21616) );
  OAI22_X2 U2099 ( .A1(n17135), .A2(n26497), .B1(n25798), .B2(n11527), .ZN(
        n21617) );
  OAI22_X2 U2100 ( .A1(n17172), .A2(n26497), .B1(n25800), .B2(n11527), .ZN(
        n21618) );
  OAI22_X2 U2101 ( .A1(n17209), .A2(n26497), .B1(n25803), .B2(n11527), .ZN(
        n21619) );
  OAI22_X2 U2102 ( .A1(n17246), .A2(n26497), .B1(n25806), .B2(n11527), .ZN(
        n21620) );
  OAI22_X2 U2103 ( .A1(n17283), .A2(n26497), .B1(n25809), .B2(n11527), .ZN(
        n21621) );
  OAI22_X2 U2104 ( .A1(n17320), .A2(n26497), .B1(n25812), .B2(n11527), .ZN(
        n21622) );
  OAI22_X2 U2105 ( .A1(n17357), .A2(n26497), .B1(n25815), .B2(n11527), .ZN(
        n21623) );
  OAI22_X2 U2106 ( .A1(n17394), .A2(n26497), .B1(n25818), .B2(n11527), .ZN(
        n21624) );
  OAI22_X2 U2107 ( .A1(n17431), .A2(n26497), .B1(n25821), .B2(n11527), .ZN(
        n21625) );
  OAI22_X2 U2108 ( .A1(n17468), .A2(n26497), .B1(n25824), .B2(n11527), .ZN(
        n21626) );
  OAI22_X2 U2109 ( .A1(n17505), .A2(n26497), .B1(n25831), .B2(n11527), .ZN(
        n21627) );
  OAI22_X2 U2110 ( .A1(n17542), .A2(n26497), .B1(n25832), .B2(n11527), .ZN(
        n21628) );
  OAI22_X2 U2113 ( .A1(n16988), .A2(n26496), .B1(n25784), .B2(n11530), .ZN(
        n21629) );
  OAI22_X2 U2114 ( .A1(n17025), .A2(n26496), .B1(n25787), .B2(n11530), .ZN(
        n21630) );
  OAI22_X2 U2115 ( .A1(n17062), .A2(n26496), .B1(n25790), .B2(n11530), .ZN(
        n21631) );
  OAI22_X2 U2116 ( .A1(n17099), .A2(n26496), .B1(n25794), .B2(n11530), .ZN(
        n21632) );
  OAI22_X2 U2117 ( .A1(n17136), .A2(n26496), .B1(n25799), .B2(n11530), .ZN(
        n21633) );
  OAI22_X2 U2118 ( .A1(n17173), .A2(n26496), .B1(n25802), .B2(n11530), .ZN(
        n21634) );
  OAI22_X2 U2119 ( .A1(n17210), .A2(n26496), .B1(n25805), .B2(n11530), .ZN(
        n21635) );
  OAI22_X2 U2120 ( .A1(n17247), .A2(n26496), .B1(n25808), .B2(n11530), .ZN(
        n21636) );
  OAI22_X2 U2121 ( .A1(n17284), .A2(n26496), .B1(n25811), .B2(n11530), .ZN(
        n21637) );
  OAI22_X2 U2122 ( .A1(n17321), .A2(n26496), .B1(n25814), .B2(n11530), .ZN(
        n21638) );
  OAI22_X2 U2123 ( .A1(n17358), .A2(n26496), .B1(n25817), .B2(n11530), .ZN(
        n21639) );
  OAI22_X2 U2124 ( .A1(n17395), .A2(n26496), .B1(n25820), .B2(n11530), .ZN(
        n21640) );
  OAI22_X2 U2125 ( .A1(n17432), .A2(n26496), .B1(n25823), .B2(n11530), .ZN(
        n21641) );
  OAI22_X2 U2126 ( .A1(n17469), .A2(n26496), .B1(n25826), .B2(n11530), .ZN(
        n21642) );
  OAI22_X2 U2127 ( .A1(n17506), .A2(n26496), .B1(n25830), .B2(n11530), .ZN(
        n21643) );
  OAI22_X2 U2128 ( .A1(n17543), .A2(n26496), .B1(n25834), .B2(n11530), .ZN(
        n21644) );
  OAI22_X2 U2131 ( .A1(n16992), .A2(n26495), .B1(n25782), .B2(n11532), .ZN(
        n21645) );
  OAI22_X2 U2132 ( .A1(n17029), .A2(n26495), .B1(n25785), .B2(n11532), .ZN(
        n21646) );
  OAI22_X2 U2133 ( .A1(n17066), .A2(n26495), .B1(n25788), .B2(n11532), .ZN(
        n21647) );
  OAI22_X2 U2134 ( .A1(n17103), .A2(n26495), .B1(n25791), .B2(n11532), .ZN(
        n21648) );
  OAI22_X2 U2135 ( .A1(n17140), .A2(n26495), .B1(n25796), .B2(n11532), .ZN(
        n21649) );
  OAI22_X2 U2136 ( .A1(n17177), .A2(n26495), .B1(n25800), .B2(n11532), .ZN(
        n21650) );
  OAI22_X2 U2137 ( .A1(n17214), .A2(n26495), .B1(n25803), .B2(n11532), .ZN(
        n21651) );
  OAI22_X2 U2138 ( .A1(n17251), .A2(n26495), .B1(n25806), .B2(n11532), .ZN(
        n21652) );
  OAI22_X2 U2139 ( .A1(n17288), .A2(n26495), .B1(n25809), .B2(n11532), .ZN(
        n21653) );
  OAI22_X2 U2140 ( .A1(n17325), .A2(n26495), .B1(n25812), .B2(n11532), .ZN(
        n21654) );
  OAI22_X2 U2141 ( .A1(n17362), .A2(n26495), .B1(n25815), .B2(n11532), .ZN(
        n21655) );
  OAI22_X2 U2142 ( .A1(n17399), .A2(n26495), .B1(n25818), .B2(n11532), .ZN(
        n21656) );
  OAI22_X2 U2143 ( .A1(n17436), .A2(n26495), .B1(n25821), .B2(n11532), .ZN(
        n21657) );
  OAI22_X2 U2144 ( .A1(n17473), .A2(n26495), .B1(n25824), .B2(n11532), .ZN(
        n21658) );
  OAI22_X2 U2145 ( .A1(n17510), .A2(n26495), .B1(n25827), .B2(n11532), .ZN(
        n21659) );
  OAI22_X2 U2146 ( .A1(n17547), .A2(n26495), .B1(n25832), .B2(n11532), .ZN(
        n21660) );
  OAI22_X2 U2149 ( .A1(n16993), .A2(n26494), .B1(n25784), .B2(n11534), .ZN(
        n21661) );
  OAI22_X2 U2150 ( .A1(n17030), .A2(n26494), .B1(n25787), .B2(n11534), .ZN(
        n21662) );
  OAI22_X2 U2151 ( .A1(n17067), .A2(n26494), .B1(n25790), .B2(n11534), .ZN(
        n21663) );
  OAI22_X2 U2152 ( .A1(n17104), .A2(n26494), .B1(n25791), .B2(n11534), .ZN(
        n21664) );
  OAI22_X2 U2153 ( .A1(n17141), .A2(n26494), .B1(n25796), .B2(n11534), .ZN(
        n21665) );
  OAI22_X2 U2154 ( .A1(n17178), .A2(n26494), .B1(n25802), .B2(n11534), .ZN(
        n21666) );
  OAI22_X2 U2155 ( .A1(n17215), .A2(n26494), .B1(n25805), .B2(n11534), .ZN(
        n21667) );
  OAI22_X2 U2156 ( .A1(n17252), .A2(n26494), .B1(n25808), .B2(n11534), .ZN(
        n21668) );
  OAI22_X2 U2157 ( .A1(n17289), .A2(n26494), .B1(n25811), .B2(n11534), .ZN(
        n21669) );
  OAI22_X2 U2158 ( .A1(n17326), .A2(n26494), .B1(n25814), .B2(n11534), .ZN(
        n21670) );
  OAI22_X2 U2159 ( .A1(n17363), .A2(n26494), .B1(n25817), .B2(n11534), .ZN(
        n21671) );
  OAI22_X2 U2160 ( .A1(n17400), .A2(n26494), .B1(n25820), .B2(n11534), .ZN(
        n21672) );
  OAI22_X2 U2161 ( .A1(n17437), .A2(n26494), .B1(n25823), .B2(n11534), .ZN(
        n21673) );
  OAI22_X2 U2162 ( .A1(n17474), .A2(n26494), .B1(n25826), .B2(n11534), .ZN(
        n21674) );
  OAI22_X2 U2163 ( .A1(n17511), .A2(n26494), .B1(n25827), .B2(n11534), .ZN(
        n21675) );
  OAI22_X2 U2164 ( .A1(n17548), .A2(n26494), .B1(n25834), .B2(n11534), .ZN(
        n21676) );
  OAI22_X2 U2167 ( .A1(n16386), .A2(n26431), .B1(n25784), .B2(n11536), .ZN(
        n21677) );
  OAI22_X2 U2168 ( .A1(n16423), .A2(n26431), .B1(n25787), .B2(n11536), .ZN(
        n21678) );
  OAI22_X2 U2169 ( .A1(n16460), .A2(n26431), .B1(n25790), .B2(n11536), .ZN(
        n21679) );
  OAI22_X2 U2170 ( .A1(n16497), .A2(n26431), .B1(n25792), .B2(n11536), .ZN(
        n21680) );
  OAI22_X2 U2171 ( .A1(n16534), .A2(n26431), .B1(n25797), .B2(n11536), .ZN(
        n21681) );
  OAI22_X2 U2172 ( .A1(n16571), .A2(n26431), .B1(n25802), .B2(n11536), .ZN(
        n21682) );
  OAI22_X2 U2173 ( .A1(n16608), .A2(n26431), .B1(n25805), .B2(n11536), .ZN(
        n21683) );
  OAI22_X2 U2174 ( .A1(n16645), .A2(n26431), .B1(n25808), .B2(n11536), .ZN(
        n21684) );
  OAI22_X2 U2175 ( .A1(n16682), .A2(n26431), .B1(n25811), .B2(n11536), .ZN(
        n21685) );
  OAI22_X2 U2176 ( .A1(n16719), .A2(n26431), .B1(n25814), .B2(n11536), .ZN(
        n21686) );
  OAI22_X2 U2177 ( .A1(n16756), .A2(n26431), .B1(n25817), .B2(n11536), .ZN(
        n21687) );
  OAI22_X2 U2178 ( .A1(n16793), .A2(n26431), .B1(n25820), .B2(n11536), .ZN(
        n21688) );
  OAI22_X2 U2179 ( .A1(n16830), .A2(n26431), .B1(n25823), .B2(n11536), .ZN(
        n21689) );
  OAI22_X2 U2180 ( .A1(n16867), .A2(n26431), .B1(n25826), .B2(n11536), .ZN(
        n21690) );
  OAI22_X2 U2181 ( .A1(n16904), .A2(n26431), .B1(n25828), .B2(n11536), .ZN(
        n21691) );
  OAI22_X2 U2182 ( .A1(n16941), .A2(n26431), .B1(n25834), .B2(n11536), .ZN(
        n21692) );
  OAI22_X2 U2185 ( .A1(n16387), .A2(n26430), .B1(n25783), .B2(n11539), .ZN(
        n21693) );
  OAI22_X2 U2186 ( .A1(n16424), .A2(n26430), .B1(n25786), .B2(n11539), .ZN(
        n21694) );
  OAI22_X2 U2187 ( .A1(n16461), .A2(n26430), .B1(n25789), .B2(n11539), .ZN(
        n21695) );
  OAI22_X2 U2188 ( .A1(n16498), .A2(n26430), .B1(n25795), .B2(n11539), .ZN(
        n21696) );
  OAI22_X2 U2189 ( .A1(n16535), .A2(n26430), .B1(n25797), .B2(n11539), .ZN(
        n21697) );
  OAI22_X2 U2190 ( .A1(n16572), .A2(n26430), .B1(n25801), .B2(n11539), .ZN(
        n21698) );
  OAI22_X2 U2191 ( .A1(n16609), .A2(n26430), .B1(n25804), .B2(n11539), .ZN(
        n21699) );
  OAI22_X2 U2192 ( .A1(n16646), .A2(n26430), .B1(n25807), .B2(n11539), .ZN(
        n21700) );
  OAI22_X2 U2193 ( .A1(n16683), .A2(n26430), .B1(n25810), .B2(n11539), .ZN(
        n21701) );
  OAI22_X2 U2194 ( .A1(n16720), .A2(n26430), .B1(n25813), .B2(n11539), .ZN(
        n21702) );
  OAI22_X2 U2195 ( .A1(n16757), .A2(n26430), .B1(n25816), .B2(n11539), .ZN(
        n21703) );
  OAI22_X2 U2196 ( .A1(n16794), .A2(n26430), .B1(n25819), .B2(n11539), .ZN(
        n21704) );
  OAI22_X2 U2197 ( .A1(n16831), .A2(n26430), .B1(n25822), .B2(n11539), .ZN(
        n21705) );
  OAI22_X2 U2198 ( .A1(n16868), .A2(n26430), .B1(n25825), .B2(n11539), .ZN(
        n21706) );
  OAI22_X2 U2199 ( .A1(n16905), .A2(n26430), .B1(n25831), .B2(n11539), .ZN(
        n21707) );
  OAI22_X2 U2200 ( .A1(n16942), .A2(n26430), .B1(n25833), .B2(n11539), .ZN(
        n21708) );
  OAI22_X2 U2203 ( .A1(n16391), .A2(n26429), .B1(n25783), .B2(n11541), .ZN(
        n21709) );
  OAI22_X2 U2204 ( .A1(n16428), .A2(n26429), .B1(n25786), .B2(n11541), .ZN(
        n21710) );
  OAI22_X2 U2205 ( .A1(n16465), .A2(n26429), .B1(n25789), .B2(n11541), .ZN(
        n21711) );
  OAI22_X2 U2206 ( .A1(n16502), .A2(n26429), .B1(n25794), .B2(n11541), .ZN(
        n21712) );
  OAI22_X2 U2207 ( .A1(n16539), .A2(n26429), .B1(n25799), .B2(n11541), .ZN(
        n21713) );
  OAI22_X2 U2208 ( .A1(n16576), .A2(n26429), .B1(n25801), .B2(n11541), .ZN(
        n21714) );
  OAI22_X2 U2209 ( .A1(n16613), .A2(n26429), .B1(n25804), .B2(n11541), .ZN(
        n21715) );
  OAI22_X2 U2210 ( .A1(n16650), .A2(n26429), .B1(n25807), .B2(n11541), .ZN(
        n21716) );
  OAI22_X2 U2211 ( .A1(n16687), .A2(n26429), .B1(n25810), .B2(n11541), .ZN(
        n21717) );
  OAI22_X2 U2212 ( .A1(n16724), .A2(n26429), .B1(n25813), .B2(n11541), .ZN(
        n21718) );
  OAI22_X2 U2213 ( .A1(n16761), .A2(n26429), .B1(n25816), .B2(n11541), .ZN(
        n21719) );
  OAI22_X2 U2214 ( .A1(n16798), .A2(n26429), .B1(n25819), .B2(n11541), .ZN(
        n21720) );
  OAI22_X2 U2215 ( .A1(n16835), .A2(n26429), .B1(n25822), .B2(n11541), .ZN(
        n21721) );
  OAI22_X2 U2216 ( .A1(n16872), .A2(n26429), .B1(n25825), .B2(n11541), .ZN(
        n21722) );
  OAI22_X2 U2217 ( .A1(n16909), .A2(n26429), .B1(n25830), .B2(n11541), .ZN(
        n21723) );
  OAI22_X2 U2218 ( .A1(n16946), .A2(n26429), .B1(n25833), .B2(n11541), .ZN(
        n21724) );
  OAI22_X2 U2221 ( .A1(n16392), .A2(n26428), .B1(n25783), .B2(n11543), .ZN(
        n21725) );
  OAI22_X2 U2222 ( .A1(n16429), .A2(n26428), .B1(n25786), .B2(n11543), .ZN(
        n21726) );
  OAI22_X2 U2223 ( .A1(n16466), .A2(n26428), .B1(n25789), .B2(n11543), .ZN(
        n21727) );
  OAI22_X2 U2224 ( .A1(n16503), .A2(n26428), .B1(n25791), .B2(n11543), .ZN(
        n21728) );
  OAI22_X2 U2225 ( .A1(n16540), .A2(n26428), .B1(n25796), .B2(n11543), .ZN(
        n21729) );
  OAI22_X2 U2226 ( .A1(n16577), .A2(n26428), .B1(n25801), .B2(n11543), .ZN(
        n21730) );
  OAI22_X2 U2227 ( .A1(n16614), .A2(n26428), .B1(n25804), .B2(n11543), .ZN(
        n21731) );
  OAI22_X2 U2228 ( .A1(n16651), .A2(n26428), .B1(n25807), .B2(n11543), .ZN(
        n21732) );
  OAI22_X2 U2229 ( .A1(n16688), .A2(n26428), .B1(n25810), .B2(n11543), .ZN(
        n21733) );
  OAI22_X2 U2230 ( .A1(n16725), .A2(n26428), .B1(n25813), .B2(n11543), .ZN(
        n21734) );
  OAI22_X2 U2231 ( .A1(n16762), .A2(n26428), .B1(n25816), .B2(n11543), .ZN(
        n21735) );
  OAI22_X2 U2232 ( .A1(n16799), .A2(n26428), .B1(n25819), .B2(n11543), .ZN(
        n21736) );
  OAI22_X2 U2233 ( .A1(n16836), .A2(n26428), .B1(n25822), .B2(n11543), .ZN(
        n21737) );
  OAI22_X2 U2234 ( .A1(n16873), .A2(n26428), .B1(n25825), .B2(n11543), .ZN(
        n21738) );
  OAI22_X2 U2235 ( .A1(n16910), .A2(n26428), .B1(n25827), .B2(n11543), .ZN(
        n21739) );
  OAI22_X2 U2236 ( .A1(n16947), .A2(n26428), .B1(n25833), .B2(n11543), .ZN(
        n21740) );
  OAI22_X2 U2239 ( .A1(n18162), .A2(n26440), .B1(n25782), .B2(n11545), .ZN(
        n21741) );
  OAI22_X2 U2240 ( .A1(n18199), .A2(n26440), .B1(n25785), .B2(n11545), .ZN(
        n21742) );
  OAI22_X2 U2241 ( .A1(n18236), .A2(n26440), .B1(n25788), .B2(n11545), .ZN(
        n21743) );
  OAI22_X2 U2242 ( .A1(n18273), .A2(n26440), .B1(n25792), .B2(n11545), .ZN(
        n21744) );
  OAI22_X2 U2243 ( .A1(n18310), .A2(n26440), .B1(n25797), .B2(n11545), .ZN(
        n21745) );
  OAI22_X2 U2244 ( .A1(n18347), .A2(n26440), .B1(n25800), .B2(n11545), .ZN(
        n21746) );
  OAI22_X2 U2245 ( .A1(n18384), .A2(n26440), .B1(n25803), .B2(n11545), .ZN(
        n21747) );
  OAI22_X2 U2246 ( .A1(n18421), .A2(n26440), .B1(n25806), .B2(n11545), .ZN(
        n21748) );
  OAI22_X2 U2247 ( .A1(n18458), .A2(n26440), .B1(n25809), .B2(n11545), .ZN(
        n21749) );
  OAI22_X2 U2248 ( .A1(n18495), .A2(n26440), .B1(n25812), .B2(n11545), .ZN(
        n21750) );
  OAI22_X2 U2249 ( .A1(n18532), .A2(n26440), .B1(n25815), .B2(n11545), .ZN(
        n21751) );
  OAI22_X2 U2250 ( .A1(n18569), .A2(n26440), .B1(n25818), .B2(n11545), .ZN(
        n21752) );
  OAI22_X2 U2251 ( .A1(n18606), .A2(n26440), .B1(n25821), .B2(n11545), .ZN(
        n21753) );
  OAI22_X2 U2252 ( .A1(n18643), .A2(n26440), .B1(n25824), .B2(n11545), .ZN(
        n21754) );
  OAI22_X2 U2253 ( .A1(n18680), .A2(n26440), .B1(n25828), .B2(n11545), .ZN(
        n21755) );
  OAI22_X2 U2254 ( .A1(n18717), .A2(n26440), .B1(n25832), .B2(n11545), .ZN(
        n21756) );
  OAI22_X2 U2257 ( .A1(n18163), .A2(n26439), .B1(n25782), .B2(n11548), .ZN(
        n21757) );
  OAI22_X2 U2258 ( .A1(n18200), .A2(n26439), .B1(n25785), .B2(n11548), .ZN(
        n21758) );
  OAI22_X2 U2259 ( .A1(n18237), .A2(n26439), .B1(n25788), .B2(n11548), .ZN(
        n21759) );
  OAI22_X2 U2260 ( .A1(n18274), .A2(n26439), .B1(n25795), .B2(n11548), .ZN(
        n21760) );
  OAI22_X2 U2261 ( .A1(n18311), .A2(n26439), .B1(n25799), .B2(n11548), .ZN(
        n21761) );
  OAI22_X2 U2262 ( .A1(n18348), .A2(n26439), .B1(n25800), .B2(n11548), .ZN(
        n21762) );
  OAI22_X2 U2263 ( .A1(n18385), .A2(n26439), .B1(n25803), .B2(n11548), .ZN(
        n21763) );
  OAI22_X2 U2264 ( .A1(n18422), .A2(n26439), .B1(n25806), .B2(n11548), .ZN(
        n21764) );
  OAI22_X2 U2265 ( .A1(n18459), .A2(n26439), .B1(n25809), .B2(n11548), .ZN(
        n21765) );
  OAI22_X2 U2266 ( .A1(n18496), .A2(n26439), .B1(n25812), .B2(n11548), .ZN(
        n21766) );
  OAI22_X2 U2267 ( .A1(n18533), .A2(n26439), .B1(n25815), .B2(n11548), .ZN(
        n21767) );
  OAI22_X2 U2268 ( .A1(n18570), .A2(n26439), .B1(n25818), .B2(n11548), .ZN(
        n21768) );
  OAI22_X2 U2269 ( .A1(n18607), .A2(n26439), .B1(n25821), .B2(n11548), .ZN(
        n21769) );
  OAI22_X2 U2270 ( .A1(n18644), .A2(n26439), .B1(n25824), .B2(n11548), .ZN(
        n21770) );
  OAI22_X2 U2271 ( .A1(n18681), .A2(n26439), .B1(n25831), .B2(n11548), .ZN(
        n21771) );
  OAI22_X2 U2272 ( .A1(n18718), .A2(n26439), .B1(n25832), .B2(n11548), .ZN(
        n21772) );
  OAI22_X2 U2275 ( .A1(n18167), .A2(n26438), .B1(n25782), .B2(n11550), .ZN(
        n21773) );
  OAI22_X2 U2276 ( .A1(n18204), .A2(n26438), .B1(n25785), .B2(n11550), .ZN(
        n21774) );
  OAI22_X2 U2277 ( .A1(n18241), .A2(n26438), .B1(n25788), .B2(n11550), .ZN(
        n21775) );
  OAI22_X2 U2278 ( .A1(n18278), .A2(n26438), .B1(n25793), .B2(n11550), .ZN(
        n21776) );
  OAI22_X2 U2279 ( .A1(n18315), .A2(n26438), .B1(n25798), .B2(n11550), .ZN(
        n21777) );
  OAI22_X2 U2280 ( .A1(n18352), .A2(n26438), .B1(n25800), .B2(n11550), .ZN(
        n21778) );
  OAI22_X2 U2281 ( .A1(n18389), .A2(n26438), .B1(n25803), .B2(n11550), .ZN(
        n21779) );
  OAI22_X2 U2282 ( .A1(n18426), .A2(n26438), .B1(n25806), .B2(n11550), .ZN(
        n21780) );
  OAI22_X2 U2283 ( .A1(n18463), .A2(n26438), .B1(n25809), .B2(n11550), .ZN(
        n21781) );
  OAI22_X2 U2284 ( .A1(n18500), .A2(n26438), .B1(n25812), .B2(n11550), .ZN(
        n21782) );
  OAI22_X2 U2285 ( .A1(n18537), .A2(n26438), .B1(n25815), .B2(n11550), .ZN(
        n21783) );
  OAI22_X2 U2286 ( .A1(n18574), .A2(n26438), .B1(n25818), .B2(n11550), .ZN(
        n21784) );
  OAI22_X2 U2287 ( .A1(n18611), .A2(n26438), .B1(n25821), .B2(n11550), .ZN(
        n21785) );
  OAI22_X2 U2288 ( .A1(n18648), .A2(n26438), .B1(n25824), .B2(n11550), .ZN(
        n21786) );
  OAI22_X2 U2289 ( .A1(n18685), .A2(n26438), .B1(n25829), .B2(n11550), .ZN(
        n21787) );
  OAI22_X2 U2290 ( .A1(n18722), .A2(n26438), .B1(n25832), .B2(n11550), .ZN(
        n21788) );
  OAI22_X2 U2293 ( .A1(n18168), .A2(n26437), .B1(n25784), .B2(n11552), .ZN(
        n21789) );
  OAI22_X2 U2294 ( .A1(n18205), .A2(n26437), .B1(n25787), .B2(n11552), .ZN(
        n21790) );
  OAI22_X2 U2295 ( .A1(n18242), .A2(n26437), .B1(n25790), .B2(n11552), .ZN(
        n21791) );
  OAI22_X2 U2296 ( .A1(n18279), .A2(n26437), .B1(n25791), .B2(n11552), .ZN(
        n21792) );
  OAI22_X2 U2297 ( .A1(n18316), .A2(n26437), .B1(n25796), .B2(n11552), .ZN(
        n21793) );
  OAI22_X2 U2298 ( .A1(n18353), .A2(n26437), .B1(n25802), .B2(n11552), .ZN(
        n21794) );
  OAI22_X2 U2299 ( .A1(n18390), .A2(n26437), .B1(n25805), .B2(n11552), .ZN(
        n21795) );
  OAI22_X2 U2300 ( .A1(n18427), .A2(n26437), .B1(n25808), .B2(n11552), .ZN(
        n21796) );
  OAI22_X2 U2301 ( .A1(n18464), .A2(n26437), .B1(n25811), .B2(n11552), .ZN(
        n21797) );
  OAI22_X2 U2302 ( .A1(n18501), .A2(n26437), .B1(n25814), .B2(n11552), .ZN(
        n21798) );
  OAI22_X2 U2303 ( .A1(n18538), .A2(n26437), .B1(n25817), .B2(n11552), .ZN(
        n21799) );
  OAI22_X2 U2304 ( .A1(n18575), .A2(n26437), .B1(n25820), .B2(n11552), .ZN(
        n21800) );
  OAI22_X2 U2305 ( .A1(n18612), .A2(n26437), .B1(n25823), .B2(n11552), .ZN(
        n21801) );
  OAI22_X2 U2306 ( .A1(n18649), .A2(n26437), .B1(n25826), .B2(n11552), .ZN(
        n21802) );
  OAI22_X2 U2307 ( .A1(n18686), .A2(n26437), .B1(n25827), .B2(n11552), .ZN(
        n21803) );
  OAI22_X2 U2308 ( .A1(n18723), .A2(n26437), .B1(n25834), .B2(n11552), .ZN(
        n21804) );
  OAI22_X2 U2311 ( .A1(n17570), .A2(n26449), .B1(n25784), .B2(n11554), .ZN(
        n21805) );
  OAI22_X2 U2312 ( .A1(n17607), .A2(n26449), .B1(n25787), .B2(n11554), .ZN(
        n21806) );
  OAI22_X2 U2313 ( .A1(n17644), .A2(n26449), .B1(n25790), .B2(n11554), .ZN(
        n21807) );
  OAI22_X2 U2314 ( .A1(n17681), .A2(n26449), .B1(n25792), .B2(n11554), .ZN(
        n21808) );
  OAI22_X2 U2315 ( .A1(n17718), .A2(n26449), .B1(n25797), .B2(n11554), .ZN(
        n21809) );
  OAI22_X2 U2316 ( .A1(n17755), .A2(n26449), .B1(n25802), .B2(n11554), .ZN(
        n21810) );
  OAI22_X2 U2317 ( .A1(n17792), .A2(n26449), .B1(n25805), .B2(n11554), .ZN(
        n21811) );
  OAI22_X2 U2318 ( .A1(n17829), .A2(n26449), .B1(n25808), .B2(n11554), .ZN(
        n21812) );
  OAI22_X2 U2319 ( .A1(n17866), .A2(n26449), .B1(n25811), .B2(n11554), .ZN(
        n21813) );
  OAI22_X2 U2320 ( .A1(n17903), .A2(n26449), .B1(n25814), .B2(n11554), .ZN(
        n21814) );
  OAI22_X2 U2321 ( .A1(n17940), .A2(n26449), .B1(n25817), .B2(n11554), .ZN(
        n21815) );
  OAI22_X2 U2322 ( .A1(n17977), .A2(n26449), .B1(n25820), .B2(n11554), .ZN(
        n21816) );
  OAI22_X2 U2323 ( .A1(n18014), .A2(n26449), .B1(n25823), .B2(n11554), .ZN(
        n21817) );
  OAI22_X2 U2324 ( .A1(n18051), .A2(n26449), .B1(n25826), .B2(n11554), .ZN(
        n21818) );
  OAI22_X2 U2325 ( .A1(n18088), .A2(n26449), .B1(n25828), .B2(n11554), .ZN(
        n21819) );
  OAI22_X2 U2326 ( .A1(n18125), .A2(n26449), .B1(n25834), .B2(n11554), .ZN(
        n21820) );
  OAI22_X2 U2329 ( .A1(n17571), .A2(n26448), .B1(n25783), .B2(n11557), .ZN(
        n21821) );
  OAI22_X2 U2330 ( .A1(n17608), .A2(n26448), .B1(n25786), .B2(n11557), .ZN(
        n21822) );
  OAI22_X2 U2331 ( .A1(n17645), .A2(n26448), .B1(n25789), .B2(n11557), .ZN(
        n21823) );
  OAI22_X2 U2332 ( .A1(n17682), .A2(n26448), .B1(n25795), .B2(n11557), .ZN(
        n21824) );
  OAI22_X2 U2333 ( .A1(n17719), .A2(n26448), .B1(n25797), .B2(n11557), .ZN(
        n21825) );
  OAI22_X2 U2334 ( .A1(n17756), .A2(n26448), .B1(n25801), .B2(n11557), .ZN(
        n21826) );
  OAI22_X2 U2335 ( .A1(n17793), .A2(n26448), .B1(n25804), .B2(n11557), .ZN(
        n21827) );
  OAI22_X2 U2336 ( .A1(n17830), .A2(n26448), .B1(n25807), .B2(n11557), .ZN(
        n21828) );
  OAI22_X2 U2337 ( .A1(n17867), .A2(n26448), .B1(n25810), .B2(n11557), .ZN(
        n21829) );
  OAI22_X2 U2338 ( .A1(n17904), .A2(n26448), .B1(n25813), .B2(n11557), .ZN(
        n21830) );
  OAI22_X2 U2339 ( .A1(n17941), .A2(n26448), .B1(n25816), .B2(n11557), .ZN(
        n21831) );
  OAI22_X2 U2340 ( .A1(n17978), .A2(n26448), .B1(n25819), .B2(n11557), .ZN(
        n21832) );
  OAI22_X2 U2341 ( .A1(n18015), .A2(n26448), .B1(n25822), .B2(n11557), .ZN(
        n21833) );
  OAI22_X2 U2342 ( .A1(n18052), .A2(n26448), .B1(n25825), .B2(n11557), .ZN(
        n21834) );
  OAI22_X2 U2343 ( .A1(n18089), .A2(n26448), .B1(n25831), .B2(n11557), .ZN(
        n21835) );
  OAI22_X2 U2344 ( .A1(n18126), .A2(n26448), .B1(n25833), .B2(n11557), .ZN(
        n21836) );
  OAI22_X2 U2347 ( .A1(n17575), .A2(n26447), .B1(n25783), .B2(n11559), .ZN(
        n21837) );
  OAI22_X2 U2348 ( .A1(n17612), .A2(n26447), .B1(n25786), .B2(n11559), .ZN(
        n21838) );
  OAI22_X2 U2349 ( .A1(n17649), .A2(n26447), .B1(n25789), .B2(n11559), .ZN(
        n21839) );
  OAI22_X2 U2350 ( .A1(n17686), .A2(n26447), .B1(n25793), .B2(n11559), .ZN(
        n21840) );
  OAI22_X2 U2351 ( .A1(n17723), .A2(n26447), .B1(n25798), .B2(n11559), .ZN(
        n21841) );
  OAI22_X2 U2352 ( .A1(n17760), .A2(n26447), .B1(n25801), .B2(n11559), .ZN(
        n21842) );
  OAI22_X2 U2353 ( .A1(n17797), .A2(n26447), .B1(n25804), .B2(n11559), .ZN(
        n21843) );
  OAI22_X2 U2354 ( .A1(n17834), .A2(n26447), .B1(n25807), .B2(n11559), .ZN(
        n21844) );
  OAI22_X2 U2355 ( .A1(n17871), .A2(n26447), .B1(n25810), .B2(n11559), .ZN(
        n21845) );
  OAI22_X2 U2356 ( .A1(n17908), .A2(n26447), .B1(n25813), .B2(n11559), .ZN(
        n21846) );
  OAI22_X2 U2357 ( .A1(n17945), .A2(n26447), .B1(n25816), .B2(n11559), .ZN(
        n21847) );
  OAI22_X2 U2358 ( .A1(n17982), .A2(n26447), .B1(n25819), .B2(n11559), .ZN(
        n21848) );
  OAI22_X2 U2359 ( .A1(n18019), .A2(n26447), .B1(n25822), .B2(n11559), .ZN(
        n21849) );
  OAI22_X2 U2360 ( .A1(n18056), .A2(n26447), .B1(n25825), .B2(n11559), .ZN(
        n21850) );
  OAI22_X2 U2361 ( .A1(n18093), .A2(n26447), .B1(n25829), .B2(n11559), .ZN(
        n21851) );
  OAI22_X2 U2362 ( .A1(n18130), .A2(n26447), .B1(n25833), .B2(n11559), .ZN(
        n21852) );
  OAI22_X2 U2365 ( .A1(n17576), .A2(n26446), .B1(n25782), .B2(n11561), .ZN(
        n21853) );
  OAI22_X2 U2366 ( .A1(n17613), .A2(n26446), .B1(n25785), .B2(n11561), .ZN(
        n21854) );
  OAI22_X2 U2367 ( .A1(n17650), .A2(n26446), .B1(n25788), .B2(n11561), .ZN(
        n21855) );
  OAI22_X2 U2368 ( .A1(n17687), .A2(n26446), .B1(n25791), .B2(n11561), .ZN(
        n21856) );
  OAI22_X2 U2369 ( .A1(n17724), .A2(n26446), .B1(n25796), .B2(n11561), .ZN(
        n21857) );
  OAI22_X2 U2370 ( .A1(n17761), .A2(n26446), .B1(n25800), .B2(n11561), .ZN(
        n21858) );
  OAI22_X2 U2371 ( .A1(n17798), .A2(n26446), .B1(n25803), .B2(n11561), .ZN(
        n21859) );
  OAI22_X2 U2372 ( .A1(n17835), .A2(n26446), .B1(n25806), .B2(n11561), .ZN(
        n21860) );
  OAI22_X2 U2373 ( .A1(n17872), .A2(n26446), .B1(n25809), .B2(n11561), .ZN(
        n21861) );
  OAI22_X2 U2374 ( .A1(n17909), .A2(n26446), .B1(n25812), .B2(n11561), .ZN(
        n21862) );
  OAI22_X2 U2375 ( .A1(n17946), .A2(n26446), .B1(n25815), .B2(n11561), .ZN(
        n21863) );
  OAI22_X2 U2376 ( .A1(n17983), .A2(n26446), .B1(n25818), .B2(n11561), .ZN(
        n21864) );
  OAI22_X2 U2377 ( .A1(n18020), .A2(n26446), .B1(n25821), .B2(n11561), .ZN(
        n21865) );
  OAI22_X2 U2378 ( .A1(n18057), .A2(n26446), .B1(n25824), .B2(n11561), .ZN(
        n21866) );
  OAI22_X2 U2379 ( .A1(n18094), .A2(n26446), .B1(n25827), .B2(n11561), .ZN(
        n21867) );
  OAI22_X2 U2380 ( .A1(n18131), .A2(n26446), .B1(n25832), .B2(n11561), .ZN(
        n21868) );
  OAI22_X2 U2383 ( .A1(n16978), .A2(n26458), .B1(n25784), .B2(n11563), .ZN(
        n21869) );
  OAI22_X2 U2384 ( .A1(n17015), .A2(n26458), .B1(n25787), .B2(n11563), .ZN(
        n21870) );
  OAI22_X2 U2385 ( .A1(n17052), .A2(n26458), .B1(n25790), .B2(n11563), .ZN(
        n21871) );
  OAI22_X2 U2386 ( .A1(n17089), .A2(n26458), .B1(n25792), .B2(n11563), .ZN(
        n21872) );
  OAI22_X2 U2387 ( .A1(n17126), .A2(n26458), .B1(n25797), .B2(n11563), .ZN(
        n21873) );
  OAI22_X2 U2388 ( .A1(n17163), .A2(n26458), .B1(n25802), .B2(n11563), .ZN(
        n21874) );
  OAI22_X2 U2389 ( .A1(n17200), .A2(n26458), .B1(n25805), .B2(n11563), .ZN(
        n21875) );
  OAI22_X2 U2390 ( .A1(n17237), .A2(n26458), .B1(n25808), .B2(n11563), .ZN(
        n21876) );
  OAI22_X2 U2391 ( .A1(n17274), .A2(n26458), .B1(n25811), .B2(n11563), .ZN(
        n21877) );
  OAI22_X2 U2392 ( .A1(n17311), .A2(n26458), .B1(n25814), .B2(n11563), .ZN(
        n21878) );
  OAI22_X2 U2393 ( .A1(n17348), .A2(n26458), .B1(n25817), .B2(n11563), .ZN(
        n21879) );
  OAI22_X2 U2394 ( .A1(n17385), .A2(n26458), .B1(n25820), .B2(n11563), .ZN(
        n21880) );
  OAI22_X2 U2395 ( .A1(n17422), .A2(n26458), .B1(n25823), .B2(n11563), .ZN(
        n21881) );
  OAI22_X2 U2396 ( .A1(n17459), .A2(n26458), .B1(n25826), .B2(n11563), .ZN(
        n21882) );
  OAI22_X2 U2397 ( .A1(n17496), .A2(n26458), .B1(n25828), .B2(n11563), .ZN(
        n21883) );
  OAI22_X2 U2398 ( .A1(n17533), .A2(n26458), .B1(n25834), .B2(n11563), .ZN(
        n21884) );
  OAI22_X2 U2401 ( .A1(n16979), .A2(n26457), .B1(n25782), .B2(n11566), .ZN(
        n21885) );
  OAI22_X2 U2402 ( .A1(n17016), .A2(n26457), .B1(n25785), .B2(n11566), .ZN(
        n21886) );
  OAI22_X2 U2403 ( .A1(n17053), .A2(n26457), .B1(n25788), .B2(n11566), .ZN(
        n21887) );
  OAI22_X2 U2404 ( .A1(n17090), .A2(n26457), .B1(n25795), .B2(n11566), .ZN(
        n21888) );
  OAI22_X2 U2405 ( .A1(n17127), .A2(n26457), .B1(n25796), .B2(n11566), .ZN(
        n21889) );
  OAI22_X2 U2406 ( .A1(n17164), .A2(n26457), .B1(n25800), .B2(n11566), .ZN(
        n21890) );
  OAI22_X2 U2407 ( .A1(n17201), .A2(n26457), .B1(n25803), .B2(n11566), .ZN(
        n21891) );
  OAI22_X2 U2408 ( .A1(n17238), .A2(n26457), .B1(n25806), .B2(n11566), .ZN(
        n21892) );
  OAI22_X2 U2409 ( .A1(n17275), .A2(n26457), .B1(n25809), .B2(n11566), .ZN(
        n21893) );
  OAI22_X2 U2410 ( .A1(n17312), .A2(n26457), .B1(n25812), .B2(n11566), .ZN(
        n21894) );
  OAI22_X2 U2411 ( .A1(n17349), .A2(n26457), .B1(n25815), .B2(n11566), .ZN(
        n21895) );
  OAI22_X2 U2412 ( .A1(n17386), .A2(n26457), .B1(n25818), .B2(n11566), .ZN(
        n21896) );
  OAI22_X2 U2413 ( .A1(n17423), .A2(n26457), .B1(n25821), .B2(n11566), .ZN(
        n21897) );
  OAI22_X2 U2414 ( .A1(n17460), .A2(n26457), .B1(n25824), .B2(n11566), .ZN(
        n21898) );
  OAI22_X2 U2415 ( .A1(n17497), .A2(n26457), .B1(n25831), .B2(n11566), .ZN(
        n21899) );
  OAI22_X2 U2416 ( .A1(n17534), .A2(n26457), .B1(n25832), .B2(n11566), .ZN(
        n21900) );
  OAI22_X2 U2419 ( .A1(n16983), .A2(n26456), .B1(n25784), .B2(n11568), .ZN(
        n21901) );
  OAI22_X2 U2420 ( .A1(n17020), .A2(n26456), .B1(n25787), .B2(n11568), .ZN(
        n21902) );
  OAI22_X2 U2421 ( .A1(n17057), .A2(n26456), .B1(n25790), .B2(n11568), .ZN(
        n21903) );
  OAI22_X2 U2422 ( .A1(n17094), .A2(n26456), .B1(n25793), .B2(n11568), .ZN(
        n21904) );
  OAI22_X2 U2423 ( .A1(n17131), .A2(n26456), .B1(n25798), .B2(n11568), .ZN(
        n21905) );
  OAI22_X2 U2424 ( .A1(n17168), .A2(n26456), .B1(n25802), .B2(n11568), .ZN(
        n21906) );
  OAI22_X2 U2425 ( .A1(n17205), .A2(n26456), .B1(n25805), .B2(n11568), .ZN(
        n21907) );
  OAI22_X2 U2426 ( .A1(n17242), .A2(n26456), .B1(n25808), .B2(n11568), .ZN(
        n21908) );
  OAI22_X2 U2427 ( .A1(n17279), .A2(n26456), .B1(n25811), .B2(n11568), .ZN(
        n21909) );
  OAI22_X2 U2428 ( .A1(n17316), .A2(n26456), .B1(n25814), .B2(n11568), .ZN(
        n21910) );
  OAI22_X2 U2429 ( .A1(n17353), .A2(n26456), .B1(n25817), .B2(n11568), .ZN(
        n21911) );
  OAI22_X2 U2430 ( .A1(n17390), .A2(n26456), .B1(n25820), .B2(n11568), .ZN(
        n21912) );
  OAI22_X2 U2431 ( .A1(n17427), .A2(n26456), .B1(n25823), .B2(n11568), .ZN(
        n21913) );
  OAI22_X2 U2432 ( .A1(n17464), .A2(n26456), .B1(n25826), .B2(n11568), .ZN(
        n21914) );
  OAI22_X2 U2433 ( .A1(n17501), .A2(n26456), .B1(n25829), .B2(n11568), .ZN(
        n21915) );
  OAI22_X2 U2434 ( .A1(n17538), .A2(n26456), .B1(n25834), .B2(n11568), .ZN(
        n21916) );
  OAI22_X2 U2437 ( .A1(n16984), .A2(n26455), .B1(n25784), .B2(n11570), .ZN(
        n21917) );
  OAI22_X2 U2438 ( .A1(n17021), .A2(n26455), .B1(n25787), .B2(n11570), .ZN(
        n21918) );
  OAI22_X2 U2439 ( .A1(n17058), .A2(n26455), .B1(n25790), .B2(n11570), .ZN(
        n21919) );
  OAI22_X2 U2440 ( .A1(n17095), .A2(n26455), .B1(n25791), .B2(n11570), .ZN(
        n21920) );
  OAI22_X2 U2441 ( .A1(n17132), .A2(n26455), .B1(n25796), .B2(n11570), .ZN(
        n21921) );
  OAI22_X2 U2442 ( .A1(n17169), .A2(n26455), .B1(n25802), .B2(n11570), .ZN(
        n21922) );
  OAI22_X2 U2443 ( .A1(n17206), .A2(n26455), .B1(n25805), .B2(n11570), .ZN(
        n21923) );
  OAI22_X2 U2444 ( .A1(n17243), .A2(n26455), .B1(n25808), .B2(n11570), .ZN(
        n21924) );
  OAI22_X2 U2445 ( .A1(n17280), .A2(n26455), .B1(n25811), .B2(n11570), .ZN(
        n21925) );
  OAI22_X2 U2446 ( .A1(n17317), .A2(n26455), .B1(n25814), .B2(n11570), .ZN(
        n21926) );
  OAI22_X2 U2447 ( .A1(n17354), .A2(n26455), .B1(n25817), .B2(n11570), .ZN(
        n21927) );
  OAI22_X2 U2448 ( .A1(n17391), .A2(n26455), .B1(n25820), .B2(n11570), .ZN(
        n21928) );
  OAI22_X2 U2449 ( .A1(n17428), .A2(n26455), .B1(n25823), .B2(n11570), .ZN(
        n21929) );
  OAI22_X2 U2450 ( .A1(n17465), .A2(n26455), .B1(n25826), .B2(n11570), .ZN(
        n21930) );
  OAI22_X2 U2451 ( .A1(n17502), .A2(n26455), .B1(n25827), .B2(n11570), .ZN(
        n21931) );
  OAI22_X2 U2452 ( .A1(n17539), .A2(n26455), .B1(n25834), .B2(n11570), .ZN(
        n21932) );
  OAI22_X2 U2455 ( .A1(n16377), .A2(n26395), .B1(n25783), .B2(n11572), .ZN(
        n21933) );
  OAI22_X2 U2456 ( .A1(n16414), .A2(n26395), .B1(n25786), .B2(n11572), .ZN(
        n21934) );
  OAI22_X2 U2457 ( .A1(n16451), .A2(n26395), .B1(n25789), .B2(n11572), .ZN(
        n21935) );
  OAI22_X2 U2458 ( .A1(n16488), .A2(n26395), .B1(n25792), .B2(n11572), .ZN(
        n21936) );
  OAI22_X2 U2459 ( .A1(n16525), .A2(n26395), .B1(n25797), .B2(n11572), .ZN(
        n21937) );
  OAI22_X2 U2460 ( .A1(n16562), .A2(n26395), .B1(n25801), .B2(n11572), .ZN(
        n21938) );
  OAI22_X2 U2461 ( .A1(n16599), .A2(n26395), .B1(n25804), .B2(n11572), .ZN(
        n21939) );
  OAI22_X2 U2462 ( .A1(n16636), .A2(n26395), .B1(n25807), .B2(n11572), .ZN(
        n21940) );
  OAI22_X2 U2463 ( .A1(n16673), .A2(n26395), .B1(n25810), .B2(n11572), .ZN(
        n21941) );
  OAI22_X2 U2464 ( .A1(n16710), .A2(n26395), .B1(n25813), .B2(n11572), .ZN(
        n21942) );
  OAI22_X2 U2465 ( .A1(n16747), .A2(n26395), .B1(n25816), .B2(n11572), .ZN(
        n21943) );
  OAI22_X2 U2466 ( .A1(n16784), .A2(n26395), .B1(n25819), .B2(n11572), .ZN(
        n21944) );
  OAI22_X2 U2467 ( .A1(n16821), .A2(n26395), .B1(n25822), .B2(n11572), .ZN(
        n21945) );
  OAI22_X2 U2468 ( .A1(n16858), .A2(n26395), .B1(n25825), .B2(n11572), .ZN(
        n21946) );
  OAI22_X2 U2469 ( .A1(n16895), .A2(n26395), .B1(n25828), .B2(n11572), .ZN(
        n21947) );
  OAI22_X2 U2470 ( .A1(n16932), .A2(n26395), .B1(n25833), .B2(n11572), .ZN(
        n21948) );
  OAI22_X2 U2473 ( .A1(n16378), .A2(n26394), .B1(n25782), .B2(n11575), .ZN(
        n21949) );
  OAI22_X2 U2474 ( .A1(n16415), .A2(n26394), .B1(n25785), .B2(n11575), .ZN(
        n21950) );
  OAI22_X2 U2475 ( .A1(n16452), .A2(n26394), .B1(n25788), .B2(n11575), .ZN(
        n21951) );
  OAI22_X2 U2476 ( .A1(n16489), .A2(n26394), .B1(n25795), .B2(n11575), .ZN(
        n21952) );
  OAI22_X2 U2477 ( .A1(n16526), .A2(n26394), .B1(n25798), .B2(n11575), .ZN(
        n21953) );
  OAI22_X2 U2478 ( .A1(n16563), .A2(n26394), .B1(n25800), .B2(n11575), .ZN(
        n21954) );
  OAI22_X2 U2479 ( .A1(n16600), .A2(n26394), .B1(n25803), .B2(n11575), .ZN(
        n21955) );
  OAI22_X2 U2480 ( .A1(n16637), .A2(n26394), .B1(n25806), .B2(n11575), .ZN(
        n21956) );
  OAI22_X2 U2481 ( .A1(n16674), .A2(n26394), .B1(n25809), .B2(n11575), .ZN(
        n21957) );
  OAI22_X2 U2482 ( .A1(n16711), .A2(n26394), .B1(n25812), .B2(n11575), .ZN(
        n21958) );
  OAI22_X2 U2483 ( .A1(n16748), .A2(n26394), .B1(n25815), .B2(n11575), .ZN(
        n21959) );
  OAI22_X2 U2484 ( .A1(n16785), .A2(n26394), .B1(n25818), .B2(n11575), .ZN(
        n21960) );
  OAI22_X2 U2485 ( .A1(n16822), .A2(n26394), .B1(n25821), .B2(n11575), .ZN(
        n21961) );
  OAI22_X2 U2486 ( .A1(n16859), .A2(n26394), .B1(n25824), .B2(n11575), .ZN(
        n21962) );
  OAI22_X2 U2487 ( .A1(n16896), .A2(n26394), .B1(n25831), .B2(n11575), .ZN(
        n21963) );
  OAI22_X2 U2488 ( .A1(n16933), .A2(n26394), .B1(n25832), .B2(n11575), .ZN(
        n21964) );
  OAI22_X2 U2491 ( .A1(n16382), .A2(n26393), .B1(n25783), .B2(n11577), .ZN(
        n21965) );
  OAI22_X2 U2492 ( .A1(n16419), .A2(n26393), .B1(n25786), .B2(n11577), .ZN(
        n21966) );
  OAI22_X2 U2493 ( .A1(n16456), .A2(n26393), .B1(n25789), .B2(n11577), .ZN(
        n21967) );
  OAI22_X2 U2494 ( .A1(n16493), .A2(n26393), .B1(n25793), .B2(n11577), .ZN(
        n21968) );
  OAI22_X2 U2495 ( .A1(n16530), .A2(n26393), .B1(n25798), .B2(n11577), .ZN(
        n21969) );
  OAI22_X2 U2496 ( .A1(n16567), .A2(n26393), .B1(n25801), .B2(n11577), .ZN(
        n21970) );
  OAI22_X2 U2497 ( .A1(n16604), .A2(n26393), .B1(n25804), .B2(n11577), .ZN(
        n21971) );
  OAI22_X2 U2498 ( .A1(n16641), .A2(n26393), .B1(n25807), .B2(n11577), .ZN(
        n21972) );
  OAI22_X2 U2499 ( .A1(n16678), .A2(n26393), .B1(n25810), .B2(n11577), .ZN(
        n21973) );
  OAI22_X2 U2500 ( .A1(n16715), .A2(n26393), .B1(n25813), .B2(n11577), .ZN(
        n21974) );
  OAI22_X2 U2501 ( .A1(n16752), .A2(n26393), .B1(n25816), .B2(n11577), .ZN(
        n21975) );
  OAI22_X2 U2502 ( .A1(n16789), .A2(n26393), .B1(n25819), .B2(n11577), .ZN(
        n21976) );
  OAI22_X2 U2503 ( .A1(n16826), .A2(n26393), .B1(n25822), .B2(n11577), .ZN(
        n21977) );
  OAI22_X2 U2504 ( .A1(n16863), .A2(n26393), .B1(n25825), .B2(n11577), .ZN(
        n21978) );
  OAI22_X2 U2505 ( .A1(n16900), .A2(n26393), .B1(n25829), .B2(n11577), .ZN(
        n21979) );
  OAI22_X2 U2506 ( .A1(n16937), .A2(n26393), .B1(n25833), .B2(n11577), .ZN(
        n21980) );
  OAI22_X2 U2509 ( .A1(n16383), .A2(n26392), .B1(n25782), .B2(n11579), .ZN(
        n21981) );
  OAI22_X2 U2510 ( .A1(n16420), .A2(n26392), .B1(n25785), .B2(n11579), .ZN(
        n21982) );
  OAI22_X2 U2511 ( .A1(n16457), .A2(n26392), .B1(n25788), .B2(n11579), .ZN(
        n21983) );
  OAI22_X2 U2512 ( .A1(n16494), .A2(n26392), .B1(n25792), .B2(n11579), .ZN(
        n21984) );
  OAI22_X2 U2513 ( .A1(n16531), .A2(n26392), .B1(n25797), .B2(n11579), .ZN(
        n21985) );
  OAI22_X2 U2514 ( .A1(n16568), .A2(n26392), .B1(n25800), .B2(n11579), .ZN(
        n21986) );
  OAI22_X2 U2515 ( .A1(n16605), .A2(n26392), .B1(n25803), .B2(n11579), .ZN(
        n21987) );
  OAI22_X2 U2516 ( .A1(n16642), .A2(n26392), .B1(n25806), .B2(n11579), .ZN(
        n21988) );
  OAI22_X2 U2517 ( .A1(n16679), .A2(n26392), .B1(n25809), .B2(n11579), .ZN(
        n21989) );
  OAI22_X2 U2518 ( .A1(n16716), .A2(n26392), .B1(n25812), .B2(n11579), .ZN(
        n21990) );
  OAI22_X2 U2519 ( .A1(n16753), .A2(n26392), .B1(n25815), .B2(n11579), .ZN(
        n21991) );
  OAI22_X2 U2520 ( .A1(n16790), .A2(n26392), .B1(n25818), .B2(n11579), .ZN(
        n21992) );
  OAI22_X2 U2521 ( .A1(n16827), .A2(n26392), .B1(n25821), .B2(n11579), .ZN(
        n21993) );
  OAI22_X2 U2522 ( .A1(n16864), .A2(n26392), .B1(n25824), .B2(n11579), .ZN(
        n21994) );
  OAI22_X2 U2523 ( .A1(n16901), .A2(n26392), .B1(n25828), .B2(n11579), .ZN(
        n21995) );
  OAI22_X2 U2524 ( .A1(n16938), .A2(n26392), .B1(n25832), .B2(n11579), .ZN(
        n21996) );
  OAI22_X2 U2527 ( .A1(n18153), .A2(n26404), .B1(n25783), .B2(n11581), .ZN(
        n21997) );
  OAI22_X2 U2528 ( .A1(n18190), .A2(n26404), .B1(n25786), .B2(n11581), .ZN(
        n21998) );
  OAI22_X2 U2529 ( .A1(n18227), .A2(n26404), .B1(n25789), .B2(n11581), .ZN(
        n21999) );
  OAI22_X2 U2530 ( .A1(n18264), .A2(n26404), .B1(n25791), .B2(n11581), .ZN(
        n22000) );
  OAI22_X2 U2531 ( .A1(n18301), .A2(n26404), .B1(n25796), .B2(n11581), .ZN(
        n22001) );
  OAI22_X2 U2532 ( .A1(n18338), .A2(n26404), .B1(n25801), .B2(n11581), .ZN(
        n22002) );
  OAI22_X2 U2533 ( .A1(n18375), .A2(n26404), .B1(n25804), .B2(n11581), .ZN(
        n22003) );
  OAI22_X2 U2534 ( .A1(n18412), .A2(n26404), .B1(n25807), .B2(n11581), .ZN(
        n22004) );
  OAI22_X2 U2535 ( .A1(n18449), .A2(n26404), .B1(n25810), .B2(n11581), .ZN(
        n22005) );
  OAI22_X2 U2536 ( .A1(n18486), .A2(n26404), .B1(n25813), .B2(n11581), .ZN(
        n22006) );
  OAI22_X2 U2537 ( .A1(n18523), .A2(n26404), .B1(n25816), .B2(n11581), .ZN(
        n22007) );
  OAI22_X2 U2538 ( .A1(n18560), .A2(n26404), .B1(n25819), .B2(n11581), .ZN(
        n22008) );
  OAI22_X2 U2539 ( .A1(n18597), .A2(n26404), .B1(n25822), .B2(n11581), .ZN(
        n22009) );
  OAI22_X2 U2540 ( .A1(n18634), .A2(n26404), .B1(n25825), .B2(n11581), .ZN(
        n22010) );
  OAI22_X2 U2541 ( .A1(n18671), .A2(n26404), .B1(n25827), .B2(n11581), .ZN(
        n22011) );
  OAI22_X2 U2542 ( .A1(n18708), .A2(n26404), .B1(n25833), .B2(n11581), .ZN(
        n22012) );
  OAI22_X2 U2545 ( .A1(n18154), .A2(n26403), .B1(n25784), .B2(n11584), .ZN(
        n22013) );
  OAI22_X2 U2546 ( .A1(n18191), .A2(n26403), .B1(n25787), .B2(n11584), .ZN(
        n22014) );
  OAI22_X2 U2547 ( .A1(n18228), .A2(n26403), .B1(n25790), .B2(n11584), .ZN(
        n22015) );
  OAI22_X2 U2548 ( .A1(n18265), .A2(n26403), .B1(n25792), .B2(n11584), .ZN(
        n22016) );
  OAI22_X2 U2549 ( .A1(n18302), .A2(n26403), .B1(n25797), .B2(n11584), .ZN(
        n22017) );
  OAI22_X2 U2550 ( .A1(n18339), .A2(n26403), .B1(n25802), .B2(n11584), .ZN(
        n22018) );
  OAI22_X2 U2551 ( .A1(n18376), .A2(n26403), .B1(n25805), .B2(n11584), .ZN(
        n22019) );
  OAI22_X2 U2552 ( .A1(n18413), .A2(n26403), .B1(n25808), .B2(n11584), .ZN(
        n22020) );
  OAI22_X2 U2553 ( .A1(n18450), .A2(n26403), .B1(n25811), .B2(n11584), .ZN(
        n22021) );
  OAI22_X2 U2554 ( .A1(n18487), .A2(n26403), .B1(n25814), .B2(n11584), .ZN(
        n22022) );
  OAI22_X2 U2555 ( .A1(n18524), .A2(n26403), .B1(n25817), .B2(n11584), .ZN(
        n22023) );
  OAI22_X2 U2556 ( .A1(n18561), .A2(n26403), .B1(n25820), .B2(n11584), .ZN(
        n22024) );
  OAI22_X2 U2557 ( .A1(n18598), .A2(n26403), .B1(n25823), .B2(n11584), .ZN(
        n22025) );
  OAI22_X2 U2558 ( .A1(n18635), .A2(n26403), .B1(n25826), .B2(n11584), .ZN(
        n22026) );
  OAI22_X2 U2559 ( .A1(n18672), .A2(n26403), .B1(n25828), .B2(n11584), .ZN(
        n22027) );
  OAI22_X2 U2560 ( .A1(n18709), .A2(n26403), .B1(n25834), .B2(n11584), .ZN(
        n22028) );
  OAI22_X2 U2563 ( .A1(n18158), .A2(n26402), .B1(n25784), .B2(n11586), .ZN(
        n22029) );
  OAI22_X2 U2564 ( .A1(n18195), .A2(n26402), .B1(n25787), .B2(n11586), .ZN(
        n22030) );
  OAI22_X2 U2565 ( .A1(n18232), .A2(n26402), .B1(n25790), .B2(n11586), .ZN(
        n22031) );
  OAI22_X2 U2566 ( .A1(n18269), .A2(n26402), .B1(n25795), .B2(n11586), .ZN(
        n22032) );
  OAI22_X2 U2567 ( .A1(n18306), .A2(n26402), .B1(n25799), .B2(n11586), .ZN(
        n22033) );
  OAI22_X2 U2568 ( .A1(n18343), .A2(n26402), .B1(n25802), .B2(n11586), .ZN(
        n22034) );
  OAI22_X2 U2569 ( .A1(n18380), .A2(n26402), .B1(n25805), .B2(n11586), .ZN(
        n22035) );
  OAI22_X2 U2570 ( .A1(n18417), .A2(n26402), .B1(n25808), .B2(n11586), .ZN(
        n22036) );
  OAI22_X2 U2571 ( .A1(n18454), .A2(n26402), .B1(n25811), .B2(n11586), .ZN(
        n22037) );
  OAI22_X2 U2572 ( .A1(n18491), .A2(n26402), .B1(n25814), .B2(n11586), .ZN(
        n22038) );
  OAI22_X2 U2573 ( .A1(n18528), .A2(n26402), .B1(n25817), .B2(n11586), .ZN(
        n22039) );
  OAI22_X2 U2574 ( .A1(n18565), .A2(n26402), .B1(n25820), .B2(n11586), .ZN(
        n22040) );
  OAI22_X2 U2575 ( .A1(n18602), .A2(n26402), .B1(n25823), .B2(n11586), .ZN(
        n22041) );
  OAI22_X2 U2576 ( .A1(n18639), .A2(n26402), .B1(n25826), .B2(n11586), .ZN(
        n22042) );
  OAI22_X2 U2577 ( .A1(n18676), .A2(n26402), .B1(n25831), .B2(n11586), .ZN(
        n22043) );
  OAI22_X2 U2578 ( .A1(n18713), .A2(n26402), .B1(n25834), .B2(n11586), .ZN(
        n22044) );
  OAI22_X2 U2581 ( .A1(n18159), .A2(n26401), .B1(n25782), .B2(n11588), .ZN(
        n22045) );
  OAI22_X2 U2582 ( .A1(n18196), .A2(n26401), .B1(n25785), .B2(n11588), .ZN(
        n22046) );
  OAI22_X2 U2583 ( .A1(n18233), .A2(n26401), .B1(n25788), .B2(n11588), .ZN(
        n22047) );
  OAI22_X2 U2584 ( .A1(n18270), .A2(n26401), .B1(n25794), .B2(n11588), .ZN(
        n22048) );
  OAI22_X2 U2585 ( .A1(n18307), .A2(n26401), .B1(n25799), .B2(n11588), .ZN(
        n22049) );
  OAI22_X2 U2586 ( .A1(n18344), .A2(n26401), .B1(n25800), .B2(n11588), .ZN(
        n22050) );
  OAI22_X2 U2587 ( .A1(n18381), .A2(n26401), .B1(n25803), .B2(n11588), .ZN(
        n22051) );
  OAI22_X2 U2588 ( .A1(n18418), .A2(n26401), .B1(n25806), .B2(n11588), .ZN(
        n22052) );
  OAI22_X2 U2589 ( .A1(n18455), .A2(n26401), .B1(n25809), .B2(n11588), .ZN(
        n22053) );
  OAI22_X2 U2590 ( .A1(n18492), .A2(n26401), .B1(n25812), .B2(n11588), .ZN(
        n22054) );
  OAI22_X2 U2591 ( .A1(n18529), .A2(n26401), .B1(n25815), .B2(n11588), .ZN(
        n22055) );
  OAI22_X2 U2592 ( .A1(n18566), .A2(n26401), .B1(n25818), .B2(n11588), .ZN(
        n22056) );
  OAI22_X2 U2593 ( .A1(n18603), .A2(n26401), .B1(n25821), .B2(n11588), .ZN(
        n22057) );
  OAI22_X2 U2594 ( .A1(n18640), .A2(n26401), .B1(n25824), .B2(n11588), .ZN(
        n22058) );
  OAI22_X2 U2595 ( .A1(n18677), .A2(n26401), .B1(n25830), .B2(n11588), .ZN(
        n22059) );
  OAI22_X2 U2596 ( .A1(n18714), .A2(n26401), .B1(n25832), .B2(n11588), .ZN(
        n22060) );
  OAI22_X2 U2599 ( .A1(n17561), .A2(n26413), .B1(n25783), .B2(n11590), .ZN(
        n22061) );
  OAI22_X2 U2600 ( .A1(n17598), .A2(n26413), .B1(n25786), .B2(n11590), .ZN(
        n22062) );
  OAI22_X2 U2601 ( .A1(n17635), .A2(n26413), .B1(n25789), .B2(n11590), .ZN(
        n22063) );
  OAI22_X2 U2602 ( .A1(n17672), .A2(n26413), .B1(n25792), .B2(n11590), .ZN(
        n22064) );
  OAI22_X2 U2603 ( .A1(n17709), .A2(n26413), .B1(n25797), .B2(n11590), .ZN(
        n22065) );
  OAI22_X2 U2604 ( .A1(n17746), .A2(n26413), .B1(n25801), .B2(n11590), .ZN(
        n22066) );
  OAI22_X2 U2605 ( .A1(n17783), .A2(n26413), .B1(n25804), .B2(n11590), .ZN(
        n22067) );
  OAI22_X2 U2606 ( .A1(n17820), .A2(n26413), .B1(n25807), .B2(n11590), .ZN(
        n22068) );
  OAI22_X2 U2607 ( .A1(n17857), .A2(n26413), .B1(n25810), .B2(n11590), .ZN(
        n22069) );
  OAI22_X2 U2608 ( .A1(n17894), .A2(n26413), .B1(n25813), .B2(n11590), .ZN(
        n22070) );
  OAI22_X2 U2609 ( .A1(n17931), .A2(n26413), .B1(n25816), .B2(n11590), .ZN(
        n22071) );
  OAI22_X2 U2610 ( .A1(n17968), .A2(n26413), .B1(n25819), .B2(n11590), .ZN(
        n22072) );
  OAI22_X2 U2611 ( .A1(n18005), .A2(n26413), .B1(n25822), .B2(n11590), .ZN(
        n22073) );
  OAI22_X2 U2612 ( .A1(n18042), .A2(n26413), .B1(n25825), .B2(n11590), .ZN(
        n22074) );
  OAI22_X2 U2613 ( .A1(n18079), .A2(n26413), .B1(n25828), .B2(n11590), .ZN(
        n22075) );
  OAI22_X2 U2614 ( .A1(n18116), .A2(n26413), .B1(n25833), .B2(n11590), .ZN(
        n22076) );
  OAI22_X2 U2617 ( .A1(n17562), .A2(n26412), .B1(n25782), .B2(n11593), .ZN(
        n22077) );
  OAI22_X2 U2618 ( .A1(n17599), .A2(n26412), .B1(n25785), .B2(n11593), .ZN(
        n22078) );
  OAI22_X2 U2619 ( .A1(n17636), .A2(n26412), .B1(n25788), .B2(n11593), .ZN(
        n22079) );
  OAI22_X2 U2620 ( .A1(n17673), .A2(n26412), .B1(n25795), .B2(n11593), .ZN(
        n22080) );
  OAI22_X2 U2621 ( .A1(n17710), .A2(n26412), .B1(n25797), .B2(n11593), .ZN(
        n22081) );
  OAI22_X2 U2622 ( .A1(n17747), .A2(n26412), .B1(n25800), .B2(n11593), .ZN(
        n22082) );
  OAI22_X2 U2623 ( .A1(n17784), .A2(n26412), .B1(n25803), .B2(n11593), .ZN(
        n22083) );
  OAI22_X2 U2624 ( .A1(n17821), .A2(n26412), .B1(n25806), .B2(n11593), .ZN(
        n22084) );
  OAI22_X2 U2625 ( .A1(n17858), .A2(n26412), .B1(n25809), .B2(n11593), .ZN(
        n22085) );
  OAI22_X2 U2626 ( .A1(n17895), .A2(n26412), .B1(n25812), .B2(n11593), .ZN(
        n22086) );
  OAI22_X2 U2627 ( .A1(n17932), .A2(n26412), .B1(n25815), .B2(n11593), .ZN(
        n22087) );
  OAI22_X2 U2628 ( .A1(n17969), .A2(n26412), .B1(n25818), .B2(n11593), .ZN(
        n22088) );
  OAI22_X2 U2629 ( .A1(n18006), .A2(n26412), .B1(n25821), .B2(n11593), .ZN(
        n22089) );
  OAI22_X2 U2630 ( .A1(n18043), .A2(n26412), .B1(n25824), .B2(n11593), .ZN(
        n22090) );
  OAI22_X2 U2631 ( .A1(n18080), .A2(n26412), .B1(n25831), .B2(n11593), .ZN(
        n22091) );
  OAI22_X2 U2632 ( .A1(n18117), .A2(n26412), .B1(n25832), .B2(n11593), .ZN(
        n22092) );
  OAI22_X2 U2635 ( .A1(n17566), .A2(n26411), .B1(n25784), .B2(n11595), .ZN(
        n22093) );
  OAI22_X2 U2636 ( .A1(n17603), .A2(n26411), .B1(n25787), .B2(n11595), .ZN(
        n22094) );
  OAI22_X2 U2637 ( .A1(n17640), .A2(n26411), .B1(n25790), .B2(n11595), .ZN(
        n22095) );
  OAI22_X2 U2638 ( .A1(n17677), .A2(n26411), .B1(n25791), .B2(n11595), .ZN(
        n22096) );
  OAI22_X2 U2639 ( .A1(n17714), .A2(n26411), .B1(n25796), .B2(n11595), .ZN(
        n22097) );
  OAI22_X2 U2640 ( .A1(n17751), .A2(n26411), .B1(n25802), .B2(n11595), .ZN(
        n22098) );
  OAI22_X2 U2641 ( .A1(n17788), .A2(n26411), .B1(n25805), .B2(n11595), .ZN(
        n22099) );
  OAI22_X2 U2642 ( .A1(n17825), .A2(n26411), .B1(n25808), .B2(n11595), .ZN(
        n22100) );
  OAI22_X2 U2643 ( .A1(n17862), .A2(n26411), .B1(n25811), .B2(n11595), .ZN(
        n22101) );
  OAI22_X2 U2644 ( .A1(n17899), .A2(n26411), .B1(n25814), .B2(n11595), .ZN(
        n22102) );
  OAI22_X2 U2645 ( .A1(n17936), .A2(n26411), .B1(n25817), .B2(n11595), .ZN(
        n22103) );
  OAI22_X2 U2646 ( .A1(n17973), .A2(n26411), .B1(n25820), .B2(n11595), .ZN(
        n22104) );
  OAI22_X2 U2647 ( .A1(n18010), .A2(n26411), .B1(n25823), .B2(n11595), .ZN(
        n22105) );
  OAI22_X2 U2648 ( .A1(n18047), .A2(n26411), .B1(n25826), .B2(n11595), .ZN(
        n22106) );
  OAI22_X2 U2649 ( .A1(n18084), .A2(n26411), .B1(n25827), .B2(n11595), .ZN(
        n22107) );
  OAI22_X2 U2650 ( .A1(n18121), .A2(n26411), .B1(n25834), .B2(n11595), .ZN(
        n22108) );
  OAI22_X2 U2653 ( .A1(n17567), .A2(n26410), .B1(n25783), .B2(n11597), .ZN(
        n22109) );
  OAI22_X2 U2654 ( .A1(n17604), .A2(n26410), .B1(n25786), .B2(n11597), .ZN(
        n22110) );
  OAI22_X2 U2655 ( .A1(n17641), .A2(n26410), .B1(n25789), .B2(n11597), .ZN(
        n22111) );
  OAI22_X2 U2656 ( .A1(n17678), .A2(n26410), .B1(n25792), .B2(n11597), .ZN(
        n22112) );
  OAI22_X2 U2657 ( .A1(n17715), .A2(n26410), .B1(n25797), .B2(n11597), .ZN(
        n22113) );
  OAI22_X2 U2658 ( .A1(n17752), .A2(n26410), .B1(n25801), .B2(n11597), .ZN(
        n22114) );
  OAI22_X2 U2659 ( .A1(n17789), .A2(n26410), .B1(n25804), .B2(n11597), .ZN(
        n22115) );
  OAI22_X2 U2660 ( .A1(n17826), .A2(n26410), .B1(n25807), .B2(n11597), .ZN(
        n22116) );
  OAI22_X2 U2661 ( .A1(n17863), .A2(n26410), .B1(n25810), .B2(n11597), .ZN(
        n22117) );
  OAI22_X2 U2662 ( .A1(n17900), .A2(n26410), .B1(n25813), .B2(n11597), .ZN(
        n22118) );
  OAI22_X2 U2663 ( .A1(n17937), .A2(n26410), .B1(n25816), .B2(n11597), .ZN(
        n22119) );
  OAI22_X2 U2664 ( .A1(n17974), .A2(n26410), .B1(n25819), .B2(n11597), .ZN(
        n22120) );
  OAI22_X2 U2665 ( .A1(n18011), .A2(n26410), .B1(n25822), .B2(n11597), .ZN(
        n22121) );
  OAI22_X2 U2666 ( .A1(n18048), .A2(n26410), .B1(n25825), .B2(n11597), .ZN(
        n22122) );
  OAI22_X2 U2667 ( .A1(n18085), .A2(n26410), .B1(n25828), .B2(n11597), .ZN(
        n22123) );
  OAI22_X2 U2668 ( .A1(n18122), .A2(n26410), .B1(n25833), .B2(n11597), .ZN(
        n22124) );
  OAI22_X2 U2671 ( .A1(n16969), .A2(n26422), .B1(n25784), .B2(n11599), .ZN(
        n22125) );
  OAI22_X2 U2672 ( .A1(n17006), .A2(n26422), .B1(n25787), .B2(n11599), .ZN(
        n22126) );
  OAI22_X2 U2673 ( .A1(n17043), .A2(n26422), .B1(n25790), .B2(n11599), .ZN(
        n22127) );
  OAI22_X2 U2674 ( .A1(n17080), .A2(n26422), .B1(n25795), .B2(n11599), .ZN(
        n22128) );
  OAI22_X2 U2675 ( .A1(n17117), .A2(n26422), .B1(n25796), .B2(n11599), .ZN(
        n22129) );
  OAI22_X2 U2676 ( .A1(n17154), .A2(n26422), .B1(n25802), .B2(n11599), .ZN(
        n22130) );
  OAI22_X2 U2677 ( .A1(n17191), .A2(n26422), .B1(n25805), .B2(n11599), .ZN(
        n22131) );
  OAI22_X2 U2678 ( .A1(n17228), .A2(n26422), .B1(n25808), .B2(n11599), .ZN(
        n22132) );
  OAI22_X2 U2679 ( .A1(n17265), .A2(n26422), .B1(n25811), .B2(n11599), .ZN(
        n22133) );
  OAI22_X2 U2680 ( .A1(n17302), .A2(n26422), .B1(n25814), .B2(n11599), .ZN(
        n22134) );
  OAI22_X2 U2681 ( .A1(n17339), .A2(n26422), .B1(n25817), .B2(n11599), .ZN(
        n22135) );
  OAI22_X2 U2682 ( .A1(n17376), .A2(n26422), .B1(n25820), .B2(n11599), .ZN(
        n22136) );
  OAI22_X2 U2683 ( .A1(n17413), .A2(n26422), .B1(n25823), .B2(n11599), .ZN(
        n22137) );
  OAI22_X2 U2684 ( .A1(n17450), .A2(n26422), .B1(n25826), .B2(n11599), .ZN(
        n22138) );
  OAI22_X2 U2685 ( .A1(n17487), .A2(n26422), .B1(n25831), .B2(n11599), .ZN(
        n22139) );
  OAI22_X2 U2686 ( .A1(n17524), .A2(n26422), .B1(n25834), .B2(n11599), .ZN(
        n22140) );
  OAI22_X2 U2689 ( .A1(n16970), .A2(n26421), .B1(n25782), .B2(n11602), .ZN(
        n22141) );
  OAI22_X2 U2690 ( .A1(n17007), .A2(n26421), .B1(n25785), .B2(n11602), .ZN(
        n22142) );
  OAI22_X2 U2691 ( .A1(n17044), .A2(n26421), .B1(n25788), .B2(n11602), .ZN(
        n22143) );
  OAI22_X2 U2692 ( .A1(n17081), .A2(n26421), .B1(n25794), .B2(n11602), .ZN(
        n22144) );
  OAI22_X2 U2693 ( .A1(n17118), .A2(n26421), .B1(n25799), .B2(n11602), .ZN(
        n22145) );
  OAI22_X2 U2694 ( .A1(n17155), .A2(n26421), .B1(n25800), .B2(n11602), .ZN(
        n22146) );
  OAI22_X2 U2695 ( .A1(n17192), .A2(n26421), .B1(n25803), .B2(n11602), .ZN(
        n22147) );
  OAI22_X2 U2696 ( .A1(n17229), .A2(n26421), .B1(n25806), .B2(n11602), .ZN(
        n22148) );
  OAI22_X2 U2697 ( .A1(n17266), .A2(n26421), .B1(n25809), .B2(n11602), .ZN(
        n22149) );
  OAI22_X2 U2698 ( .A1(n17303), .A2(n26421), .B1(n25812), .B2(n11602), .ZN(
        n22150) );
  OAI22_X2 U2699 ( .A1(n17340), .A2(n26421), .B1(n25815), .B2(n11602), .ZN(
        n22151) );
  OAI22_X2 U2700 ( .A1(n17377), .A2(n26421), .B1(n25818), .B2(n11602), .ZN(
        n22152) );
  OAI22_X2 U2701 ( .A1(n17414), .A2(n26421), .B1(n25821), .B2(n11602), .ZN(
        n22153) );
  OAI22_X2 U2702 ( .A1(n17451), .A2(n26421), .B1(n25824), .B2(n11602), .ZN(
        n22154) );
  OAI22_X2 U2703 ( .A1(n17488), .A2(n26421), .B1(n25830), .B2(n11602), .ZN(
        n22155) );
  OAI22_X2 U2704 ( .A1(n17525), .A2(n26421), .B1(n25832), .B2(n11602), .ZN(
        n22156) );
  OAI22_X2 U2707 ( .A1(n16974), .A2(n26420), .B1(n25783), .B2(n11604), .ZN(
        n22157) );
  OAI22_X2 U2708 ( .A1(n17011), .A2(n26420), .B1(n25786), .B2(n11604), .ZN(
        n22158) );
  OAI22_X2 U2709 ( .A1(n17048), .A2(n26420), .B1(n25789), .B2(n11604), .ZN(
        n22159) );
  OAI22_X2 U2710 ( .A1(n17085), .A2(n26420), .B1(n25795), .B2(n11604), .ZN(
        n22160) );
  OAI22_X2 U2711 ( .A1(n17122), .A2(n26420), .B1(n25798), .B2(n11604), .ZN(
        n22161) );
  OAI22_X2 U2712 ( .A1(n17159), .A2(n26420), .B1(n25801), .B2(n11604), .ZN(
        n22162) );
  OAI22_X2 U2713 ( .A1(n17196), .A2(n26420), .B1(n25804), .B2(n11604), .ZN(
        n22163) );
  OAI22_X2 U2714 ( .A1(n17233), .A2(n26420), .B1(n25807), .B2(n11604), .ZN(
        n22164) );
  OAI22_X2 U2715 ( .A1(n17270), .A2(n26420), .B1(n25810), .B2(n11604), .ZN(
        n22165) );
  OAI22_X2 U2716 ( .A1(n17307), .A2(n26420), .B1(n25813), .B2(n11604), .ZN(
        n22166) );
  OAI22_X2 U2717 ( .A1(n17344), .A2(n26420), .B1(n25816), .B2(n11604), .ZN(
        n22167) );
  OAI22_X2 U2718 ( .A1(n17381), .A2(n26420), .B1(n25819), .B2(n11604), .ZN(
        n22168) );
  OAI22_X2 U2719 ( .A1(n17418), .A2(n26420), .B1(n25822), .B2(n11604), .ZN(
        n22169) );
  OAI22_X2 U2720 ( .A1(n17455), .A2(n26420), .B1(n25825), .B2(n11604), .ZN(
        n22170) );
  OAI22_X2 U2721 ( .A1(n17492), .A2(n26420), .B1(n25831), .B2(n11604), .ZN(
        n22171) );
  OAI22_X2 U2722 ( .A1(n17529), .A2(n26420), .B1(n25833), .B2(n11604), .ZN(
        n22172) );
  OAI22_X2 U2725 ( .A1(n16975), .A2(n26419), .B1(n25783), .B2(n11606), .ZN(
        n22173) );
  OAI22_X2 U2726 ( .A1(n17012), .A2(n26419), .B1(n25786), .B2(n11606), .ZN(
        n22174) );
  OAI22_X2 U2727 ( .A1(n17049), .A2(n26419), .B1(n25789), .B2(n11606), .ZN(
        n22175) );
  OAI22_X2 U2728 ( .A1(n17086), .A2(n26419), .B1(n25793), .B2(n11606), .ZN(
        n22176) );
  OAI22_X2 U2729 ( .A1(n17123), .A2(n26419), .B1(n25798), .B2(n11606), .ZN(
        n22177) );
  OAI22_X2 U2730 ( .A1(n17160), .A2(n26419), .B1(n25801), .B2(n11606), .ZN(
        n22178) );
  OAI22_X2 U2731 ( .A1(n17197), .A2(n26419), .B1(n25804), .B2(n11606), .ZN(
        n22179) );
  OAI22_X2 U2732 ( .A1(n17234), .A2(n26419), .B1(n25807), .B2(n11606), .ZN(
        n22180) );
  OAI22_X2 U2733 ( .A1(n17271), .A2(n26419), .B1(n25810), .B2(n11606), .ZN(
        n22181) );
  OAI22_X2 U2734 ( .A1(n17308), .A2(n26419), .B1(n25813), .B2(n11606), .ZN(
        n22182) );
  OAI22_X2 U2735 ( .A1(n17345), .A2(n26419), .B1(n25816), .B2(n11606), .ZN(
        n22183) );
  OAI22_X2 U2736 ( .A1(n17382), .A2(n26419), .B1(n25819), .B2(n11606), .ZN(
        n22184) );
  OAI22_X2 U2737 ( .A1(n17419), .A2(n26419), .B1(n25822), .B2(n11606), .ZN(
        n22185) );
  OAI22_X2 U2738 ( .A1(n17456), .A2(n26419), .B1(n25825), .B2(n11606), .ZN(
        n22186) );
  OAI22_X2 U2739 ( .A1(n17493), .A2(n26419), .B1(n25829), .B2(n11606), .ZN(
        n22187) );
  OAI22_X2 U2740 ( .A1(n17530), .A2(n26419), .B1(n25833), .B2(n11606), .ZN(
        n22188) );
  OAI22_X2 U2743 ( .A1(n18180), .A2(n26368), .B1(n25782), .B2(n11608), .ZN(
        n22189) );
  OAI22_X2 U2744 ( .A1(n18217), .A2(n26368), .B1(n25785), .B2(n11608), .ZN(
        n22190) );
  OAI22_X2 U2745 ( .A1(n18254), .A2(n26368), .B1(n25788), .B2(n11608), .ZN(
        n22191) );
  OAI22_X2 U2746 ( .A1(n18291), .A2(n26368), .B1(n25791), .B2(n11608), .ZN(
        n22192) );
  OAI22_X2 U2747 ( .A1(n18328), .A2(n26368), .B1(n25796), .B2(n11608), .ZN(
        n22193) );
  OAI22_X2 U2748 ( .A1(n18365), .A2(n26368), .B1(n25800), .B2(n11608), .ZN(
        n22194) );
  OAI22_X2 U2749 ( .A1(n18402), .A2(n26368), .B1(n25803), .B2(n11608), .ZN(
        n22195) );
  OAI22_X2 U2750 ( .A1(n18439), .A2(n26368), .B1(n25806), .B2(n11608), .ZN(
        n22196) );
  OAI22_X2 U2751 ( .A1(n18476), .A2(n26368), .B1(n25809), .B2(n11608), .ZN(
        n22197) );
  OAI22_X2 U2752 ( .A1(n18513), .A2(n26368), .B1(n25812), .B2(n11608), .ZN(
        n22198) );
  OAI22_X2 U2753 ( .A1(n18550), .A2(n26368), .B1(n25815), .B2(n11608), .ZN(
        n22199) );
  OAI22_X2 U2754 ( .A1(n18587), .A2(n26368), .B1(n25818), .B2(n11608), .ZN(
        n22200) );
  OAI22_X2 U2755 ( .A1(n18624), .A2(n26368), .B1(n25821), .B2(n11608), .ZN(
        n22201) );
  OAI22_X2 U2756 ( .A1(n18661), .A2(n26368), .B1(n25824), .B2(n11608), .ZN(
        n22202) );
  OAI22_X2 U2757 ( .A1(n18698), .A2(n26368), .B1(n25827), .B2(n11608), .ZN(
        n22203) );
  OAI22_X2 U2758 ( .A1(n18735), .A2(n26368), .B1(n25832), .B2(n11608), .ZN(
        n22204) );
  OAI22_X2 U2761 ( .A1(n18181), .A2(n26367), .B1(n25784), .B2(n11611), .ZN(
        n22205) );
  OAI22_X2 U2762 ( .A1(n18218), .A2(n26367), .B1(n25787), .B2(n11611), .ZN(
        n22206) );
  OAI22_X2 U2763 ( .A1(n18255), .A2(n26367), .B1(n25790), .B2(n11611), .ZN(
        n22207) );
  OAI22_X2 U2764 ( .A1(n18292), .A2(n26367), .B1(n25791), .B2(n11611), .ZN(
        n22208) );
  OAI22_X2 U2765 ( .A1(n18329), .A2(n26367), .B1(n25796), .B2(n11611), .ZN(
        n22209) );
  OAI22_X2 U2766 ( .A1(n18366), .A2(n26367), .B1(n25802), .B2(n11611), .ZN(
        n22210) );
  OAI22_X2 U2767 ( .A1(n18403), .A2(n26367), .B1(n25805), .B2(n11611), .ZN(
        n22211) );
  OAI22_X2 U2768 ( .A1(n18440), .A2(n26367), .B1(n25808), .B2(n11611), .ZN(
        n22212) );
  OAI22_X2 U2769 ( .A1(n18477), .A2(n26367), .B1(n25811), .B2(n11611), .ZN(
        n22213) );
  OAI22_X2 U2770 ( .A1(n18514), .A2(n26367), .B1(n25814), .B2(n11611), .ZN(
        n22214) );
  OAI22_X2 U2771 ( .A1(n18551), .A2(n26367), .B1(n25817), .B2(n11611), .ZN(
        n22215) );
  OAI22_X2 U2772 ( .A1(n18588), .A2(n26367), .B1(n25820), .B2(n11611), .ZN(
        n22216) );
  OAI22_X2 U2773 ( .A1(n18625), .A2(n26367), .B1(n25823), .B2(n11611), .ZN(
        n22217) );
  OAI22_X2 U2774 ( .A1(n18662), .A2(n26367), .B1(n25826), .B2(n11611), .ZN(
        n22218) );
  OAI22_X2 U2775 ( .A1(n18699), .A2(n26367), .B1(n25827), .B2(n11611), .ZN(
        n22219) );
  OAI22_X2 U2776 ( .A1(n18736), .A2(n26367), .B1(n25834), .B2(n11611), .ZN(
        n22220) );
  OAI22_X2 U2779 ( .A1(n18185), .A2(n26366), .B1(n25783), .B2(n11613), .ZN(
        n22221) );
  OAI22_X2 U2780 ( .A1(n18222), .A2(n26366), .B1(n25786), .B2(n11613), .ZN(
        n22222) );
  OAI22_X2 U2781 ( .A1(n18259), .A2(n26366), .B1(n25789), .B2(n11613), .ZN(
        n22223) );
  OAI22_X2 U2782 ( .A1(n18296), .A2(n26366), .B1(n25791), .B2(n11613), .ZN(
        n22224) );
  OAI22_X2 U2783 ( .A1(n18333), .A2(n26366), .B1(n25796), .B2(n11613), .ZN(
        n22225) );
  OAI22_X2 U2784 ( .A1(n18370), .A2(n26366), .B1(n25801), .B2(n11613), .ZN(
        n22226) );
  OAI22_X2 U2785 ( .A1(n18407), .A2(n26366), .B1(n25804), .B2(n11613), .ZN(
        n22227) );
  OAI22_X2 U2786 ( .A1(n18444), .A2(n26366), .B1(n25807), .B2(n11613), .ZN(
        n22228) );
  OAI22_X2 U2787 ( .A1(n18481), .A2(n26366), .B1(n25810), .B2(n11613), .ZN(
        n22229) );
  OAI22_X2 U2788 ( .A1(n18518), .A2(n26366), .B1(n25813), .B2(n11613), .ZN(
        n22230) );
  OAI22_X2 U2789 ( .A1(n18555), .A2(n26366), .B1(n25816), .B2(n11613), .ZN(
        n22231) );
  OAI22_X2 U2790 ( .A1(n18592), .A2(n26366), .B1(n25819), .B2(n11613), .ZN(
        n22232) );
  OAI22_X2 U2791 ( .A1(n18629), .A2(n26366), .B1(n25822), .B2(n11613), .ZN(
        n22233) );
  OAI22_X2 U2792 ( .A1(n18666), .A2(n26366), .B1(n25825), .B2(n11613), .ZN(
        n22234) );
  OAI22_X2 U2793 ( .A1(n18703), .A2(n26366), .B1(n25827), .B2(n11613), .ZN(
        n22235) );
  OAI22_X2 U2794 ( .A1(n18740), .A2(n26366), .B1(n25833), .B2(n11613), .ZN(
        n22236) );
  OAI22_X2 U2797 ( .A1(n18186), .A2(n26365), .B1(n25782), .B2(n11615), .ZN(
        n22237) );
  OAI22_X2 U2798 ( .A1(n18223), .A2(n26365), .B1(n25785), .B2(n11615), .ZN(
        n22238) );
  OAI22_X2 U2799 ( .A1(n18260), .A2(n26365), .B1(n25788), .B2(n11615), .ZN(
        n22239) );
  OAI22_X2 U2800 ( .A1(n18297), .A2(n26365), .B1(n25791), .B2(n11615), .ZN(
        n22240) );
  OAI22_X2 U2801 ( .A1(n18334), .A2(n26365), .B1(n25796), .B2(n11615), .ZN(
        n22241) );
  OAI22_X2 U2802 ( .A1(n18371), .A2(n26365), .B1(n25800), .B2(n11615), .ZN(
        n22242) );
  OAI22_X2 U2803 ( .A1(n18408), .A2(n26365), .B1(n25803), .B2(n11615), .ZN(
        n22243) );
  OAI22_X2 U2804 ( .A1(n18445), .A2(n26365), .B1(n25806), .B2(n11615), .ZN(
        n22244) );
  OAI22_X2 U2805 ( .A1(n18482), .A2(n26365), .B1(n25809), .B2(n11615), .ZN(
        n22245) );
  OAI22_X2 U2806 ( .A1(n18519), .A2(n26365), .B1(n25812), .B2(n11615), .ZN(
        n22246) );
  OAI22_X2 U2807 ( .A1(n18556), .A2(n26365), .B1(n25815), .B2(n11615), .ZN(
        n22247) );
  OAI22_X2 U2808 ( .A1(n18593), .A2(n26365), .B1(n25818), .B2(n11615), .ZN(
        n22248) );
  OAI22_X2 U2809 ( .A1(n18630), .A2(n26365), .B1(n25821), .B2(n11615), .ZN(
        n22249) );
  OAI22_X2 U2810 ( .A1(n18667), .A2(n26365), .B1(n25824), .B2(n11615), .ZN(
        n22250) );
  OAI22_X2 U2811 ( .A1(n18704), .A2(n26365), .B1(n25827), .B2(n11615), .ZN(
        n22251) );
  OAI22_X2 U2812 ( .A1(n18741), .A2(n26365), .B1(n25832), .B2(n11615), .ZN(
        n22252) );
  OAI22_X2 U2815 ( .A1(n17588), .A2(n26377), .B1(n25784), .B2(n11617), .ZN(
        n22253) );
  OAI22_X2 U2816 ( .A1(n17625), .A2(n26377), .B1(n25787), .B2(n11617), .ZN(
        n22254) );
  OAI22_X2 U2817 ( .A1(n17662), .A2(n26377), .B1(n25790), .B2(n11617), .ZN(
        n22255) );
  OAI22_X2 U2818 ( .A1(n17699), .A2(n26377), .B1(n25791), .B2(n11617), .ZN(
        n22256) );
  OAI22_X2 U2819 ( .A1(n17736), .A2(n26377), .B1(n25796), .B2(n11617), .ZN(
        n22257) );
  OAI22_X2 U2820 ( .A1(n17773), .A2(n26377), .B1(n25802), .B2(n11617), .ZN(
        n22258) );
  OAI22_X2 U2821 ( .A1(n17810), .A2(n26377), .B1(n25805), .B2(n11617), .ZN(
        n22259) );
  OAI22_X2 U2822 ( .A1(n17847), .A2(n26377), .B1(n25808), .B2(n11617), .ZN(
        n22260) );
  OAI22_X2 U2823 ( .A1(n17884), .A2(n26377), .B1(n25811), .B2(n11617), .ZN(
        n22261) );
  OAI22_X2 U2824 ( .A1(n17921), .A2(n26377), .B1(n25814), .B2(n11617), .ZN(
        n22262) );
  OAI22_X2 U2825 ( .A1(n17958), .A2(n26377), .B1(n25817), .B2(n11617), .ZN(
        n22263) );
  OAI22_X2 U2826 ( .A1(n17995), .A2(n26377), .B1(n25820), .B2(n11617), .ZN(
        n22264) );
  OAI22_X2 U2827 ( .A1(n18032), .A2(n26377), .B1(n25823), .B2(n11617), .ZN(
        n22265) );
  OAI22_X2 U2828 ( .A1(n18069), .A2(n26377), .B1(n25826), .B2(n11617), .ZN(
        n22266) );
  OAI22_X2 U2829 ( .A1(n18106), .A2(n26377), .B1(n25827), .B2(n11617), .ZN(
        n22267) );
  OAI22_X2 U2830 ( .A1(n18143), .A2(n26377), .B1(n25834), .B2(n11617), .ZN(
        n22268) );
  OAI22_X2 U2833 ( .A1(n17589), .A2(n26376), .B1(n25782), .B2(n11620), .ZN(
        n22269) );
  OAI22_X2 U2834 ( .A1(n17626), .A2(n26376), .B1(n25785), .B2(n11620), .ZN(
        n22270) );
  OAI22_X2 U2835 ( .A1(n17663), .A2(n26376), .B1(n25788), .B2(n11620), .ZN(
        n22271) );
  OAI22_X2 U2836 ( .A1(n17700), .A2(n26376), .B1(n25791), .B2(n11620), .ZN(
        n22272) );
  OAI22_X2 U2837 ( .A1(n17737), .A2(n26376), .B1(n25796), .B2(n11620), .ZN(
        n22273) );
  OAI22_X2 U2838 ( .A1(n17774), .A2(n26376), .B1(n25800), .B2(n11620), .ZN(
        n22274) );
  OAI22_X2 U2839 ( .A1(n17811), .A2(n26376), .B1(n25803), .B2(n11620), .ZN(
        n22275) );
  OAI22_X2 U2840 ( .A1(n17848), .A2(n26376), .B1(n25806), .B2(n11620), .ZN(
        n22276) );
  OAI22_X2 U2841 ( .A1(n17885), .A2(n26376), .B1(n25809), .B2(n11620), .ZN(
        n22277) );
  OAI22_X2 U2842 ( .A1(n17922), .A2(n26376), .B1(n25812), .B2(n11620), .ZN(
        n22278) );
  OAI22_X2 U2843 ( .A1(n17959), .A2(n26376), .B1(n25815), .B2(n11620), .ZN(
        n22279) );
  OAI22_X2 U2844 ( .A1(n17996), .A2(n26376), .B1(n25818), .B2(n11620), .ZN(
        n22280) );
  OAI22_X2 U2845 ( .A1(n18033), .A2(n26376), .B1(n25821), .B2(n11620), .ZN(
        n22281) );
  OAI22_X2 U2846 ( .A1(n18070), .A2(n26376), .B1(n25824), .B2(n11620), .ZN(
        n22282) );
  OAI22_X2 U2847 ( .A1(n18107), .A2(n26376), .B1(n25827), .B2(n11620), .ZN(
        n22283) );
  OAI22_X2 U2848 ( .A1(n18144), .A2(n26376), .B1(n25832), .B2(n11620), .ZN(
        n22284) );
  OAI22_X2 U2851 ( .A1(n17593), .A2(n26375), .B1(n25784), .B2(n11622), .ZN(
        n22285) );
  OAI22_X2 U2852 ( .A1(n17630), .A2(n26375), .B1(n25787), .B2(n11622), .ZN(
        n22286) );
  OAI22_X2 U2853 ( .A1(n17667), .A2(n26375), .B1(n25790), .B2(n11622), .ZN(
        n22287) );
  OAI22_X2 U2854 ( .A1(n17704), .A2(n26375), .B1(n25791), .B2(n11622), .ZN(
        n22288) );
  OAI22_X2 U2855 ( .A1(n17741), .A2(n26375), .B1(n25796), .B2(n11622), .ZN(
        n22289) );
  OAI22_X2 U2856 ( .A1(n17778), .A2(n26375), .B1(n25802), .B2(n11622), .ZN(
        n22290) );
  OAI22_X2 U2857 ( .A1(n17815), .A2(n26375), .B1(n25805), .B2(n11622), .ZN(
        n22291) );
  OAI22_X2 U2858 ( .A1(n17852), .A2(n26375), .B1(n25808), .B2(n11622), .ZN(
        n22292) );
  OAI22_X2 U2859 ( .A1(n17889), .A2(n26375), .B1(n25811), .B2(n11622), .ZN(
        n22293) );
  OAI22_X2 U2860 ( .A1(n17926), .A2(n26375), .B1(n25814), .B2(n11622), .ZN(
        n22294) );
  OAI22_X2 U2861 ( .A1(n17963), .A2(n26375), .B1(n25817), .B2(n11622), .ZN(
        n22295) );
  OAI22_X2 U2862 ( .A1(n18000), .A2(n26375), .B1(n25820), .B2(n11622), .ZN(
        n22296) );
  OAI22_X2 U2863 ( .A1(n18037), .A2(n26375), .B1(n25823), .B2(n11622), .ZN(
        n22297) );
  OAI22_X2 U2864 ( .A1(n18074), .A2(n26375), .B1(n25826), .B2(n11622), .ZN(
        n22298) );
  OAI22_X2 U2865 ( .A1(n18111), .A2(n26375), .B1(n25827), .B2(n11622), .ZN(
        n22299) );
  OAI22_X2 U2866 ( .A1(n18148), .A2(n26375), .B1(n25834), .B2(n11622), .ZN(
        n22300) );
  OAI22_X2 U2869 ( .A1(n17594), .A2(n26374), .B1(n25783), .B2(n11624), .ZN(
        n22301) );
  OAI22_X2 U2870 ( .A1(n17631), .A2(n26374), .B1(n25786), .B2(n11624), .ZN(
        n22302) );
  OAI22_X2 U2871 ( .A1(n17668), .A2(n26374), .B1(n25789), .B2(n11624), .ZN(
        n22303) );
  OAI22_X2 U2872 ( .A1(n17705), .A2(n26374), .B1(n25791), .B2(n11624), .ZN(
        n22304) );
  OAI22_X2 U2873 ( .A1(n17742), .A2(n26374), .B1(n25796), .B2(n11624), .ZN(
        n22305) );
  OAI22_X2 U2874 ( .A1(n17779), .A2(n26374), .B1(n25801), .B2(n11624), .ZN(
        n22306) );
  OAI22_X2 U2875 ( .A1(n17816), .A2(n26374), .B1(n25804), .B2(n11624), .ZN(
        n22307) );
  OAI22_X2 U2876 ( .A1(n17853), .A2(n26374), .B1(n25807), .B2(n11624), .ZN(
        n22308) );
  OAI22_X2 U2877 ( .A1(n17890), .A2(n26374), .B1(n25810), .B2(n11624), .ZN(
        n22309) );
  OAI22_X2 U2878 ( .A1(n17927), .A2(n26374), .B1(n25813), .B2(n11624), .ZN(
        n22310) );
  OAI22_X2 U2879 ( .A1(n17964), .A2(n26374), .B1(n25816), .B2(n11624), .ZN(
        n22311) );
  OAI22_X2 U2880 ( .A1(n18001), .A2(n26374), .B1(n25819), .B2(n11624), .ZN(
        n22312) );
  OAI22_X2 U2881 ( .A1(n18038), .A2(n26374), .B1(n25822), .B2(n11624), .ZN(
        n22313) );
  OAI22_X2 U2882 ( .A1(n18075), .A2(n26374), .B1(n25825), .B2(n11624), .ZN(
        n22314) );
  OAI22_X2 U2883 ( .A1(n18112), .A2(n26374), .B1(n25827), .B2(n11624), .ZN(
        n22315) );
  OAI22_X2 U2884 ( .A1(n18149), .A2(n26374), .B1(n25833), .B2(n11624), .ZN(
        n22316) );
  OAI22_X2 U2887 ( .A1(n16996), .A2(n26386), .B1(n25782), .B2(n11626), .ZN(
        n22317) );
  OAI22_X2 U2888 ( .A1(n17033), .A2(n26386), .B1(n25785), .B2(n11626), .ZN(
        n22318) );
  OAI22_X2 U2889 ( .A1(n17070), .A2(n26386), .B1(n25788), .B2(n11626), .ZN(
        n22319) );
  OAI22_X2 U2890 ( .A1(n17107), .A2(n26386), .B1(n25791), .B2(n11626), .ZN(
        n22320) );
  OAI22_X2 U2891 ( .A1(n17144), .A2(n26386), .B1(n25796), .B2(n11626), .ZN(
        n22321) );
  OAI22_X2 U2892 ( .A1(n17181), .A2(n26386), .B1(n25800), .B2(n11626), .ZN(
        n22322) );
  OAI22_X2 U2893 ( .A1(n17218), .A2(n26386), .B1(n25803), .B2(n11626), .ZN(
        n22323) );
  OAI22_X2 U2894 ( .A1(n17255), .A2(n26386), .B1(n25806), .B2(n11626), .ZN(
        n22324) );
  OAI22_X2 U2895 ( .A1(n17292), .A2(n26386), .B1(n25809), .B2(n11626), .ZN(
        n22325) );
  OAI22_X2 U2896 ( .A1(n17329), .A2(n26386), .B1(n25812), .B2(n11626), .ZN(
        n22326) );
  OAI22_X2 U2897 ( .A1(n17366), .A2(n26386), .B1(n25815), .B2(n11626), .ZN(
        n22327) );
  OAI22_X2 U2898 ( .A1(n17403), .A2(n26386), .B1(n25818), .B2(n11626), .ZN(
        n22328) );
  OAI22_X2 U2899 ( .A1(n17440), .A2(n26386), .B1(n25821), .B2(n11626), .ZN(
        n22329) );
  OAI22_X2 U2900 ( .A1(n17477), .A2(n26386), .B1(n25824), .B2(n11626), .ZN(
        n22330) );
  OAI22_X2 U2901 ( .A1(n17514), .A2(n26386), .B1(n25827), .B2(n11626), .ZN(
        n22331) );
  OAI22_X2 U2902 ( .A1(n17551), .A2(n26386), .B1(n25832), .B2(n11626), .ZN(
        n22332) );
  OAI22_X2 U2905 ( .A1(n16997), .A2(n26385), .B1(n25784), .B2(n11629), .ZN(
        n22333) );
  OAI22_X2 U2906 ( .A1(n17034), .A2(n26385), .B1(n25787), .B2(n11629), .ZN(
        n22334) );
  OAI22_X2 U2907 ( .A1(n17071), .A2(n26385), .B1(n25790), .B2(n11629), .ZN(
        n22335) );
  OAI22_X2 U2908 ( .A1(n17108), .A2(n26385), .B1(n25791), .B2(n11629), .ZN(
        n22336) );
  OAI22_X2 U2909 ( .A1(n17145), .A2(n26385), .B1(n25796), .B2(n11629), .ZN(
        n22337) );
  OAI22_X2 U2910 ( .A1(n17182), .A2(n26385), .B1(n25802), .B2(n11629), .ZN(
        n22338) );
  OAI22_X2 U2911 ( .A1(n17219), .A2(n26385), .B1(n25805), .B2(n11629), .ZN(
        n22339) );
  OAI22_X2 U2912 ( .A1(n17256), .A2(n26385), .B1(n25808), .B2(n11629), .ZN(
        n22340) );
  OAI22_X2 U2913 ( .A1(n17293), .A2(n26385), .B1(n25811), .B2(n11629), .ZN(
        n22341) );
  OAI22_X2 U2914 ( .A1(n17330), .A2(n26385), .B1(n25814), .B2(n11629), .ZN(
        n22342) );
  OAI22_X2 U2915 ( .A1(n17367), .A2(n26385), .B1(n25817), .B2(n11629), .ZN(
        n22343) );
  OAI22_X2 U2916 ( .A1(n17404), .A2(n26385), .B1(n25820), .B2(n11629), .ZN(
        n22344) );
  OAI22_X2 U2917 ( .A1(n17441), .A2(n26385), .B1(n25823), .B2(n11629), .ZN(
        n22345) );
  OAI22_X2 U2918 ( .A1(n17478), .A2(n26385), .B1(n25826), .B2(n11629), .ZN(
        n22346) );
  OAI22_X2 U2919 ( .A1(n17515), .A2(n26385), .B1(n25827), .B2(n11629), .ZN(
        n22347) );
  OAI22_X2 U2920 ( .A1(n17552), .A2(n26385), .B1(n25834), .B2(n11629), .ZN(
        n22348) );
  OAI22_X2 U2923 ( .A1(n17001), .A2(n26384), .B1(n25784), .B2(n11631), .ZN(
        n22349) );
  OAI22_X2 U2924 ( .A1(n17038), .A2(n26384), .B1(n25787), .B2(n11631), .ZN(
        n22350) );
  OAI22_X2 U2925 ( .A1(n17075), .A2(n26384), .B1(n25790), .B2(n11631), .ZN(
        n22351) );
  OAI22_X2 U2926 ( .A1(n17112), .A2(n26384), .B1(n25791), .B2(n11631), .ZN(
        n22352) );
  OAI22_X2 U2927 ( .A1(n17149), .A2(n26384), .B1(n25796), .B2(n11631), .ZN(
        n22353) );
  OAI22_X2 U2928 ( .A1(n17186), .A2(n26384), .B1(n25802), .B2(n11631), .ZN(
        n22354) );
  OAI22_X2 U2929 ( .A1(n17223), .A2(n26384), .B1(n25805), .B2(n11631), .ZN(
        n22355) );
  OAI22_X2 U2930 ( .A1(n17260), .A2(n26384), .B1(n25808), .B2(n11631), .ZN(
        n22356) );
  OAI22_X2 U2931 ( .A1(n17297), .A2(n26384), .B1(n25811), .B2(n11631), .ZN(
        n22357) );
  OAI22_X2 U2932 ( .A1(n17334), .A2(n26384), .B1(n25814), .B2(n11631), .ZN(
        n22358) );
  OAI22_X2 U2933 ( .A1(n17371), .A2(n26384), .B1(n25817), .B2(n11631), .ZN(
        n22359) );
  OAI22_X2 U2934 ( .A1(n17408), .A2(n26384), .B1(n25820), .B2(n11631), .ZN(
        n22360) );
  OAI22_X2 U2935 ( .A1(n17445), .A2(n26384), .B1(n25823), .B2(n11631), .ZN(
        n22361) );
  OAI22_X2 U2936 ( .A1(n17482), .A2(n26384), .B1(n25826), .B2(n11631), .ZN(
        n22362) );
  OAI22_X2 U2937 ( .A1(n17519), .A2(n26384), .B1(n25827), .B2(n11631), .ZN(
        n22363) );
  OAI22_X2 U2938 ( .A1(n17556), .A2(n26384), .B1(n25834), .B2(n11631), .ZN(
        n22364) );
  OAI22_X2 U2941 ( .A1(n17002), .A2(n26383), .B1(n25783), .B2(n11633), .ZN(
        n22365) );
  OAI22_X2 U2942 ( .A1(n17039), .A2(n26383), .B1(n25786), .B2(n11633), .ZN(
        n22366) );
  OAI22_X2 U2943 ( .A1(n17076), .A2(n26383), .B1(n25789), .B2(n11633), .ZN(
        n22367) );
  OAI22_X2 U2944 ( .A1(n17113), .A2(n26383), .B1(n25791), .B2(n11633), .ZN(
        n22368) );
  OAI22_X2 U2945 ( .A1(n17150), .A2(n26383), .B1(n25796), .B2(n11633), .ZN(
        n22369) );
  OAI22_X2 U2946 ( .A1(n17187), .A2(n26383), .B1(n25801), .B2(n11633), .ZN(
        n22370) );
  OAI22_X2 U2947 ( .A1(n17224), .A2(n26383), .B1(n25804), .B2(n11633), .ZN(
        n22371) );
  OAI22_X2 U2948 ( .A1(n17261), .A2(n26383), .B1(n25807), .B2(n11633), .ZN(
        n22372) );
  OAI22_X2 U2949 ( .A1(n17298), .A2(n26383), .B1(n25810), .B2(n11633), .ZN(
        n22373) );
  OAI22_X2 U2950 ( .A1(n17335), .A2(n26383), .B1(n25813), .B2(n11633), .ZN(
        n22374) );
  OAI22_X2 U2951 ( .A1(n17372), .A2(n26383), .B1(n25816), .B2(n11633), .ZN(
        n22375) );
  OAI22_X2 U2952 ( .A1(n17409), .A2(n26383), .B1(n25819), .B2(n11633), .ZN(
        n22376) );
  OAI22_X2 U2953 ( .A1(n17446), .A2(n26383), .B1(n25822), .B2(n11633), .ZN(
        n22377) );
  OAI22_X2 U2954 ( .A1(n17483), .A2(n26383), .B1(n25825), .B2(n11633), .ZN(
        n22378) );
  OAI22_X2 U2955 ( .A1(n17520), .A2(n26383), .B1(n25827), .B2(n11633), .ZN(
        n22379) );
  OAI22_X2 U2956 ( .A1(n17557), .A2(n26383), .B1(n25833), .B2(n11633), .ZN(
        n22380) );
  OAI22_X2 U2960 ( .A1(n19482), .A2(n11435), .B1(n22424), .B2(n26303), .ZN(
        n22428) );
  OAI22_X2 U2961 ( .A1(n19481), .A2(n11435), .B1(n22423), .B2(n26303), .ZN(
        n22429) );
  OAI22_X2 U2962 ( .A1(n19480), .A2(n11435), .B1(n22422), .B2(n26303), .ZN(
        n22430) );
  NAND2_X2 U2963 ( .A1(n11636), .A2(n11637), .ZN(n22431) );
  AOI221_X2 U2964 ( .B1(n19476), .B2(n11638), .C1(n19475), .C2(n11639), .A(
        n11640), .ZN(n11637) );
  OAI22_X2 U2967 ( .A1(n11649), .A2(n28698), .B1(n11651), .B2(n28699), .ZN(
        n11648) );
  NAND2_X2 U2968 ( .A1(n11653), .A2(n11654), .ZN(n22432) );
  AOI221_X2 U2969 ( .B1(n19468), .B2(n11638), .C1(n19467), .C2(n11639), .A(
        n11655), .ZN(n11654) );
  OAI22_X2 U2972 ( .A1(n11649), .A2(n28706), .B1(n11651), .B2(n28707), .ZN(
        n11659) );
  NAND2_X2 U2973 ( .A1(n11662), .A2(n11663), .ZN(n22433) );
  AOI221_X2 U2974 ( .B1(n19460), .B2(n11638), .C1(n19459), .C2(n11639), .A(
        n11664), .ZN(n11663) );
  OAI22_X2 U2977 ( .A1(n11649), .A2(n28714), .B1(n11651), .B2(n28715), .ZN(
        n11668) );
  NAND2_X2 U2978 ( .A1(n11671), .A2(n11672), .ZN(n22434) );
  AOI221_X2 U2979 ( .B1(n19452), .B2(n11638), .C1(n19451), .C2(n11639), .A(
        n11673), .ZN(n11672) );
  OAI22_X2 U2982 ( .A1(n11649), .A2(n28722), .B1(n11651), .B2(n28723), .ZN(
        n11677) );
  NAND2_X2 U2983 ( .A1(n11680), .A2(n11681), .ZN(n22435) );
  AOI221_X2 U2984 ( .B1(n19444), .B2(n11638), .C1(n19443), .C2(n11639), .A(
        n11682), .ZN(n11681) );
  OAI22_X2 U2987 ( .A1(n11649), .A2(n28730), .B1(n11651), .B2(n28731), .ZN(
        n11686) );
  NAND2_X2 U2988 ( .A1(n11689), .A2(n11690), .ZN(n22436) );
  AOI221_X2 U2989 ( .B1(n19436), .B2(n11638), .C1(n19435), .C2(n11639), .A(
        n11691), .ZN(n11690) );
  OAI22_X2 U2992 ( .A1(n11649), .A2(n28738), .B1(n11651), .B2(n28739), .ZN(
        n11695) );
  NAND2_X2 U2993 ( .A1(n11698), .A2(n11699), .ZN(n22437) );
  AOI221_X2 U2994 ( .B1(n19428), .B2(n11638), .C1(n19427), .C2(n11639), .A(
        n11700), .ZN(n11699) );
  OAI22_X2 U2997 ( .A1(n11649), .A2(n28746), .B1(n11651), .B2(n28747), .ZN(
        n11704) );
  NAND2_X2 U2998 ( .A1(n11707), .A2(n11708), .ZN(n22438) );
  AOI221_X2 U2999 ( .B1(n19420), .B2(n11638), .C1(n19419), .C2(n11639), .A(
        n11709), .ZN(n11708) );
  OAI22_X2 U3002 ( .A1(n11649), .A2(n28754), .B1(n11651), .B2(n28755), .ZN(
        n11713) );
  NAND2_X2 U3003 ( .A1(n11716), .A2(n11717), .ZN(n22439) );
  AOI221_X2 U3004 ( .B1(n19412), .B2(n11638), .C1(n19411), .C2(n11639), .A(
        n11718), .ZN(n11717) );
  OAI22_X2 U3007 ( .A1(n11649), .A2(n28762), .B1(n11651), .B2(n28763), .ZN(
        n11722) );
  NAND2_X2 U3008 ( .A1(n11725), .A2(n11726), .ZN(n22440) );
  AOI221_X2 U3009 ( .B1(n19404), .B2(n11638), .C1(n19403), .C2(n11639), .A(
        n11727), .ZN(n11726) );
  OAI22_X2 U3012 ( .A1(n11649), .A2(n28770), .B1(n11651), .B2(n28771), .ZN(
        n11731) );
  NAND2_X2 U3013 ( .A1(n11734), .A2(n11735), .ZN(n22441) );
  AOI221_X2 U3014 ( .B1(n19396), .B2(n11638), .C1(n19395), .C2(n11639), .A(
        n11736), .ZN(n11735) );
  OAI22_X2 U3017 ( .A1(n11649), .A2(n28778), .B1(n11651), .B2(n28779), .ZN(
        n11740) );
  NAND2_X2 U3018 ( .A1(n11743), .A2(n11744), .ZN(n22442) );
  AOI221_X2 U3019 ( .B1(n19388), .B2(n11638), .C1(n19387), .C2(n11639), .A(
        n11745), .ZN(n11744) );
  OAI22_X2 U3022 ( .A1(n11649), .A2(n28786), .B1(n11651), .B2(n28787), .ZN(
        n11749) );
  NAND2_X2 U3023 ( .A1(n11752), .A2(n11753), .ZN(n22443) );
  AOI221_X2 U3024 ( .B1(n19380), .B2(n11638), .C1(n19379), .C2(n11639), .A(
        n11754), .ZN(n11753) );
  OAI22_X2 U3027 ( .A1(n11649), .A2(n28794), .B1(n11651), .B2(n28795), .ZN(
        n11758) );
  NAND2_X2 U3028 ( .A1(n11761), .A2(n11762), .ZN(n22444) );
  AOI221_X2 U3029 ( .B1(n19372), .B2(n11638), .C1(n19371), .C2(n11639), .A(
        n11763), .ZN(n11762) );
  OAI22_X2 U3032 ( .A1(n11649), .A2(n28802), .B1(n11651), .B2(n28803), .ZN(
        n11767) );
  NAND2_X2 U3033 ( .A1(n11770), .A2(n11771), .ZN(n22445) );
  AOI221_X2 U3034 ( .B1(n19364), .B2(n11638), .C1(n19363), .C2(n11639), .A(
        n11772), .ZN(n11771) );
  OAI22_X2 U3037 ( .A1(n11649), .A2(n28810), .B1(n11651), .B2(n28811), .ZN(
        n11776) );
  NAND2_X2 U3038 ( .A1(n11779), .A2(n11780), .ZN(n22446) );
  AOI221_X2 U3039 ( .B1(n19356), .B2(n11638), .C1(n19355), .C2(n11639), .A(
        n11781), .ZN(n11780) );
  NOR3_X2 U3043 ( .A1(n24891), .A2(n24868), .A3(n25248), .ZN(n11436) );
  OAI22_X2 U3048 ( .A1(n11649), .A2(n28817), .B1(n11651), .B2(n28818), .ZN(
        n11789) );
  NAND2_X2 U3055 ( .A1(n11283), .A2(n11793), .ZN(n22447) );
  OAI22_X2 U3074 ( .A1(n26343), .A2(n26222), .B1(n11798), .B2(n28809), .ZN(
        n22456) );
  OAI22_X2 U3076 ( .A1(n26349), .A2(n28810), .B1(n11801), .B2(n26222), .ZN(
        n22457) );
  OAI22_X2 U3078 ( .A1(n26342), .A2(n28811), .B1(n11803), .B2(n26222), .ZN(
        n22458) );
  OAI22_X2 U3080 ( .A1(n26348), .A2(n28812), .B1(n11806), .B2(n26222), .ZN(
        n22459) );
  OAI22_X2 U3082 ( .A1(n26347), .A2(n28813), .B1(n11809), .B2(n26222), .ZN(
        n22460) );
  OAI22_X2 U3084 ( .A1(n26346), .A2(n28814), .B1(n11811), .B2(n26222), .ZN(
        n22461) );
  OAI22_X2 U3086 ( .A1(n26345), .A2(n28815), .B1(n11813), .B2(n26222), .ZN(
        n22462) );
  OAI22_X2 U3088 ( .A1(n26344), .A2(n28816), .B1(n11815), .B2(n26222), .ZN(
        n22463) );
  OAI22_X2 U3091 ( .A1(n26343), .A2(n26223), .B1(n11798), .B2(n28801), .ZN(
        n22464) );
  OAI22_X2 U3093 ( .A1(n26349), .A2(n28802), .B1(n11801), .B2(n26223), .ZN(
        n22465) );
  OAI22_X2 U3095 ( .A1(n26342), .A2(n28803), .B1(n11803), .B2(n26223), .ZN(
        n22466) );
  OAI22_X2 U3097 ( .A1(n26348), .A2(n28804), .B1(n11806), .B2(n26223), .ZN(
        n22467) );
  OAI22_X2 U3099 ( .A1(n26347), .A2(n28805), .B1(n11809), .B2(n26223), .ZN(
        n22468) );
  OAI22_X2 U3101 ( .A1(n26346), .A2(n28806), .B1(n11811), .B2(n26223), .ZN(
        n22469) );
  OAI22_X2 U3103 ( .A1(n26345), .A2(n28807), .B1(n11813), .B2(n26223), .ZN(
        n22470) );
  OAI22_X2 U3105 ( .A1(n26344), .A2(n28808), .B1(n11815), .B2(n26223), .ZN(
        n22471) );
  OAI22_X2 U3108 ( .A1(n26343), .A2(n26224), .B1(n11798), .B2(n28793), .ZN(
        n22472) );
  OAI22_X2 U3110 ( .A1(n26349), .A2(n28794), .B1(n11801), .B2(n26224), .ZN(
        n22473) );
  OAI22_X2 U3112 ( .A1(n26342), .A2(n28795), .B1(n11803), .B2(n26224), .ZN(
        n22474) );
  OAI22_X2 U3114 ( .A1(n26348), .A2(n28796), .B1(n11806), .B2(n26224), .ZN(
        n22475) );
  OAI22_X2 U3116 ( .A1(n26347), .A2(n28797), .B1(n11809), .B2(n26224), .ZN(
        n22476) );
  OAI22_X2 U3118 ( .A1(n26346), .A2(n28798), .B1(n11811), .B2(n26224), .ZN(
        n22477) );
  OAI22_X2 U3120 ( .A1(n26345), .A2(n28799), .B1(n11813), .B2(n26224), .ZN(
        n22478) );
  OAI22_X2 U3122 ( .A1(n26344), .A2(n28800), .B1(n11815), .B2(n26224), .ZN(
        n22479) );
  OAI22_X2 U3125 ( .A1(n26343), .A2(n26225), .B1(n11798), .B2(n28785), .ZN(
        n22480) );
  OAI22_X2 U3127 ( .A1(n26349), .A2(n28786), .B1(n11801), .B2(n26225), .ZN(
        n22481) );
  OAI22_X2 U3129 ( .A1(n26342), .A2(n28787), .B1(n11803), .B2(n26225), .ZN(
        n22482) );
  OAI22_X2 U3131 ( .A1(n26348), .A2(n28788), .B1(n11806), .B2(n26225), .ZN(
        n22483) );
  OAI22_X2 U3133 ( .A1(n26347), .A2(n28789), .B1(n11809), .B2(n26225), .ZN(
        n22484) );
  OAI22_X2 U3135 ( .A1(n26346), .A2(n28790), .B1(n11811), .B2(n26225), .ZN(
        n22485) );
  OAI22_X2 U3137 ( .A1(n26345), .A2(n28791), .B1(n11813), .B2(n26225), .ZN(
        n22486) );
  OAI22_X2 U3139 ( .A1(n26344), .A2(n28792), .B1(n11815), .B2(n26225), .ZN(
        n22487) );
  OAI22_X2 U3142 ( .A1(n26343), .A2(n26226), .B1(n11798), .B2(n28777), .ZN(
        n22488) );
  OAI22_X2 U3144 ( .A1(n26349), .A2(n28778), .B1(n11801), .B2(n26226), .ZN(
        n22489) );
  OAI22_X2 U3146 ( .A1(n26342), .A2(n28779), .B1(n11803), .B2(n26226), .ZN(
        n22490) );
  OAI22_X2 U3148 ( .A1(n26348), .A2(n28780), .B1(n11806), .B2(n26226), .ZN(
        n22491) );
  OAI22_X2 U3150 ( .A1(n26347), .A2(n28781), .B1(n11809), .B2(n26226), .ZN(
        n22492) );
  OAI22_X2 U3152 ( .A1(n26346), .A2(n28782), .B1(n11811), .B2(n26226), .ZN(
        n22493) );
  OAI22_X2 U3154 ( .A1(n26345), .A2(n28783), .B1(n11813), .B2(n26226), .ZN(
        n22494) );
  OAI22_X2 U3156 ( .A1(n26344), .A2(n28784), .B1(n11815), .B2(n26226), .ZN(
        n22495) );
  OAI22_X2 U3159 ( .A1(n26343), .A2(n26227), .B1(n11798), .B2(n28769), .ZN(
        n22496) );
  OAI22_X2 U3161 ( .A1(n26349), .A2(n28770), .B1(n11801), .B2(n26227), .ZN(
        n22497) );
  OAI22_X2 U3163 ( .A1(n26342), .A2(n28771), .B1(n11803), .B2(n26227), .ZN(
        n22498) );
  OAI22_X2 U3165 ( .A1(n26348), .A2(n28772), .B1(n11806), .B2(n26227), .ZN(
        n22499) );
  OAI22_X2 U3167 ( .A1(n26347), .A2(n28773), .B1(n11809), .B2(n26227), .ZN(
        n22500) );
  OAI22_X2 U3169 ( .A1(n26346), .A2(n28774), .B1(n11811), .B2(n26227), .ZN(
        n22501) );
  OAI22_X2 U3171 ( .A1(n26345), .A2(n28775), .B1(n11813), .B2(n26227), .ZN(
        n22502) );
  OAI22_X2 U3173 ( .A1(n26344), .A2(n28776), .B1(n11815), .B2(n26227), .ZN(
        n22503) );
  OAI22_X2 U3176 ( .A1(n26343), .A2(n26228), .B1(n11798), .B2(n28761), .ZN(
        n22504) );
  OAI22_X2 U3178 ( .A1(n26349), .A2(n28762), .B1(n11801), .B2(n26228), .ZN(
        n22505) );
  OAI22_X2 U3180 ( .A1(n26342), .A2(n28763), .B1(n11803), .B2(n26228), .ZN(
        n22506) );
  OAI22_X2 U3182 ( .A1(n26348), .A2(n28764), .B1(n11806), .B2(n26228), .ZN(
        n22507) );
  OAI22_X2 U3184 ( .A1(n26347), .A2(n28765), .B1(n11809), .B2(n26228), .ZN(
        n22508) );
  OAI22_X2 U3186 ( .A1(n26346), .A2(n28766), .B1(n11811), .B2(n26228), .ZN(
        n22509) );
  OAI22_X2 U3188 ( .A1(n26345), .A2(n28767), .B1(n11813), .B2(n26228), .ZN(
        n22510) );
  OAI22_X2 U3190 ( .A1(n26344), .A2(n28768), .B1(n11815), .B2(n26228), .ZN(
        n22511) );
  OAI22_X2 U3193 ( .A1(n26343), .A2(n26229), .B1(n11798), .B2(n28753), .ZN(
        n22512) );
  OAI22_X2 U3195 ( .A1(n26349), .A2(n28754), .B1(n11801), .B2(n26229), .ZN(
        n22513) );
  OAI22_X2 U3197 ( .A1(n26342), .A2(n28755), .B1(n11803), .B2(n26229), .ZN(
        n22514) );
  OAI22_X2 U3199 ( .A1(n26348), .A2(n28756), .B1(n11806), .B2(n26229), .ZN(
        n22515) );
  OAI22_X2 U3201 ( .A1(n26347), .A2(n28757), .B1(n11809), .B2(n26229), .ZN(
        n22516) );
  OAI22_X2 U3203 ( .A1(n26346), .A2(n28758), .B1(n11811), .B2(n26229), .ZN(
        n22517) );
  OAI22_X2 U3205 ( .A1(n26345), .A2(n28759), .B1(n11813), .B2(n26229), .ZN(
        n22518) );
  OAI22_X2 U3207 ( .A1(n26344), .A2(n28760), .B1(n11815), .B2(n26229), .ZN(
        n22519) );
  OAI22_X2 U3210 ( .A1(n26343), .A2(n26230), .B1(n11798), .B2(n28745), .ZN(
        n22520) );
  OAI22_X2 U3212 ( .A1(n26349), .A2(n28746), .B1(n11801), .B2(n26230), .ZN(
        n22521) );
  OAI22_X2 U3214 ( .A1(n26342), .A2(n28747), .B1(n11803), .B2(n26230), .ZN(
        n22522) );
  OAI22_X2 U3216 ( .A1(n26348), .A2(n28748), .B1(n11806), .B2(n26230), .ZN(
        n22523) );
  OAI22_X2 U3218 ( .A1(n26347), .A2(n28749), .B1(n11809), .B2(n26230), .ZN(
        n22524) );
  OAI22_X2 U3220 ( .A1(n26346), .A2(n28750), .B1(n11811), .B2(n26230), .ZN(
        n22525) );
  OAI22_X2 U3222 ( .A1(n26345), .A2(n28751), .B1(n11813), .B2(n26230), .ZN(
        n22526) );
  OAI22_X2 U3224 ( .A1(n26344), .A2(n28752), .B1(n11815), .B2(n26230), .ZN(
        n22527) );
  OAI22_X2 U3227 ( .A1(n26343), .A2(n26231), .B1(n11798), .B2(n28737), .ZN(
        n22528) );
  OAI22_X2 U3229 ( .A1(n26349), .A2(n28738), .B1(n11801), .B2(n26231), .ZN(
        n22529) );
  OAI22_X2 U3231 ( .A1(n26342), .A2(n28739), .B1(n11803), .B2(n26231), .ZN(
        n22530) );
  OAI22_X2 U3233 ( .A1(n26348), .A2(n28740), .B1(n11806), .B2(n26231), .ZN(
        n22531) );
  OAI22_X2 U3235 ( .A1(n26347), .A2(n28741), .B1(n11809), .B2(n26231), .ZN(
        n22532) );
  OAI22_X2 U3237 ( .A1(n26346), .A2(n28742), .B1(n11811), .B2(n26231), .ZN(
        n22533) );
  OAI22_X2 U3239 ( .A1(n26345), .A2(n28743), .B1(n11813), .B2(n26231), .ZN(
        n22534) );
  OAI22_X2 U3241 ( .A1(n26344), .A2(n28744), .B1(n11815), .B2(n26231), .ZN(
        n22535) );
  OAI22_X2 U3244 ( .A1(n26343), .A2(n26232), .B1(n11798), .B2(n28729), .ZN(
        n22536) );
  OAI22_X2 U3246 ( .A1(n26349), .A2(n28730), .B1(n11801), .B2(n26232), .ZN(
        n22537) );
  OAI22_X2 U3248 ( .A1(n26342), .A2(n28731), .B1(n11803), .B2(n26232), .ZN(
        n22538) );
  OAI22_X2 U3250 ( .A1(n26348), .A2(n28732), .B1(n11806), .B2(n26232), .ZN(
        n22539) );
  OAI22_X2 U3252 ( .A1(n26347), .A2(n28733), .B1(n11809), .B2(n26232), .ZN(
        n22540) );
  OAI22_X2 U3254 ( .A1(n26346), .A2(n28734), .B1(n11811), .B2(n26232), .ZN(
        n22541) );
  OAI22_X2 U3256 ( .A1(n26345), .A2(n28735), .B1(n11813), .B2(n26232), .ZN(
        n22542) );
  OAI22_X2 U3258 ( .A1(n26344), .A2(n28736), .B1(n11815), .B2(n26232), .ZN(
        n22543) );
  OAI22_X2 U3261 ( .A1(n26343), .A2(n26233), .B1(n11798), .B2(n28721), .ZN(
        n22544) );
  OAI22_X2 U3263 ( .A1(n26349), .A2(n28722), .B1(n11801), .B2(n26233), .ZN(
        n22545) );
  OAI22_X2 U3265 ( .A1(n26342), .A2(n28723), .B1(n11803), .B2(n26233), .ZN(
        n22546) );
  OAI22_X2 U3267 ( .A1(n26348), .A2(n28724), .B1(n11806), .B2(n26233), .ZN(
        n22547) );
  OAI22_X2 U3269 ( .A1(n26347), .A2(n28725), .B1(n11809), .B2(n26233), .ZN(
        n22548) );
  OAI22_X2 U3271 ( .A1(n26346), .A2(n28726), .B1(n11811), .B2(n26233), .ZN(
        n22549) );
  OAI22_X2 U3273 ( .A1(n26345), .A2(n28727), .B1(n11813), .B2(n26233), .ZN(
        n22550) );
  OAI22_X2 U3275 ( .A1(n26344), .A2(n28728), .B1(n11815), .B2(n26233), .ZN(
        n22551) );
  OAI22_X2 U3278 ( .A1(n26343), .A2(n26234), .B1(n11798), .B2(n28713), .ZN(
        n22552) );
  OAI22_X2 U3280 ( .A1(n26349), .A2(n28714), .B1(n11801), .B2(n26234), .ZN(
        n22553) );
  OAI22_X2 U3282 ( .A1(n26342), .A2(n28715), .B1(n11803), .B2(n26234), .ZN(
        n22554) );
  OAI22_X2 U3284 ( .A1(n26348), .A2(n28716), .B1(n11806), .B2(n26234), .ZN(
        n22555) );
  OAI22_X2 U3286 ( .A1(n26347), .A2(n28717), .B1(n11809), .B2(n26234), .ZN(
        n22556) );
  OAI22_X2 U3288 ( .A1(n26346), .A2(n28718), .B1(n11811), .B2(n26234), .ZN(
        n22557) );
  OAI22_X2 U3290 ( .A1(n26345), .A2(n28719), .B1(n11813), .B2(n26234), .ZN(
        n22558) );
  OAI22_X2 U3292 ( .A1(n26344), .A2(n28720), .B1(n11815), .B2(n26234), .ZN(
        n22559) );
  OAI22_X2 U3295 ( .A1(n26343), .A2(n26235), .B1(n11798), .B2(n28705), .ZN(
        n22560) );
  OAI22_X2 U3297 ( .A1(n26349), .A2(n28706), .B1(n11801), .B2(n26235), .ZN(
        n22561) );
  OAI22_X2 U3299 ( .A1(n26342), .A2(n28707), .B1(n11803), .B2(n26235), .ZN(
        n22562) );
  OAI22_X2 U3301 ( .A1(n26348), .A2(n28708), .B1(n11806), .B2(n26235), .ZN(
        n22563) );
  OAI22_X2 U3303 ( .A1(n26347), .A2(n28709), .B1(n11809), .B2(n26235), .ZN(
        n22564) );
  OAI22_X2 U3305 ( .A1(n26346), .A2(n28710), .B1(n11811), .B2(n26235), .ZN(
        n22565) );
  OAI22_X2 U3307 ( .A1(n26345), .A2(n28711), .B1(n11813), .B2(n26235), .ZN(
        n22566) );
  OAI22_X2 U3309 ( .A1(n26344), .A2(n28712), .B1(n11815), .B2(n26235), .ZN(
        n22567) );
  OAI22_X2 U3312 ( .A1(n26343), .A2(n26236), .B1(n11798), .B2(n28697), .ZN(
        n22568) );
  OAI22_X2 U3314 ( .A1(n26349), .A2(n28698), .B1(n11801), .B2(n26236), .ZN(
        n22569) );
  OAI22_X2 U3318 ( .A1(n26342), .A2(n28699), .B1(n11803), .B2(n26236), .ZN(
        n22570) );
  NAND3_X2 U3321 ( .A1(n11876), .A2(n25959), .A3(n22421), .ZN(n11803) );
  OAI22_X2 U3322 ( .A1(n26348), .A2(n28700), .B1(n11806), .B2(n26236), .ZN(
        n22571) );
  NOR4_X2 U3326 ( .A1(n11878), .A2(n25958), .A3(n22420), .A4(n19348), .ZN(
        n11874) );
  OAI22_X2 U3327 ( .A1(n26347), .A2(n28701), .B1(n11809), .B2(n26236), .ZN(
        n22572) );
  OAI22_X2 U3331 ( .A1(n26346), .A2(n28702), .B1(n11811), .B2(n26236), .ZN(
        n22573) );
  NAND3_X2 U3334 ( .A1(n24894), .A2(n26129), .A3(n11880), .ZN(n11811) );
  OAI22_X2 U3335 ( .A1(n26345), .A2(n28703), .B1(n11813), .B2(n26236), .ZN(
        n22574) );
  OAI22_X2 U3339 ( .A1(n26344), .A2(n28704), .B1(n11815), .B2(n26236), .ZN(
        n22575) );
  NAND3_X2 U3343 ( .A1(n22421), .A2(n26129), .A3(n11880), .ZN(n11815) );
  NOR3_X2 U3344 ( .A1(n11878), .A2(n25958), .A3(n25255), .ZN(n11880) );
  OAI22_X2 U3370 ( .A1(n25917), .A2(n28250), .B1(n26252), .B2(n25916), .ZN(
        n22588) );
  OAI22_X2 U3372 ( .A1(n25938), .A2(n28251), .B1(n26252), .B2(n24841), .ZN(
        n22589) );
  OAI22_X2 U3374 ( .A1(n25950), .A2(n28252), .B1(n26252), .B2(n25949), .ZN(
        n22590) );
  OAI22_X2 U3376 ( .A1(n24846), .A2(n26252), .B1(n25956), .B2(n28253), .ZN(
        n22591) );
  OAI22_X2 U3387 ( .A1(n25917), .A2(n28242), .B1(n26253), .B2(n25916), .ZN(
        n22596) );
  OAI22_X2 U3389 ( .A1(n25938), .A2(n28243), .B1(n26253), .B2(n24841), .ZN(
        n22597) );
  OAI22_X2 U3393 ( .A1(n25955), .A2(n26253), .B1(n25956), .B2(n28245), .ZN(
        n22599) );
  OAI22_X2 U3396 ( .A1(n25926), .A2(n28230), .B1(n26254), .B2(n24838), .ZN(
        n22600) );
  OAI22_X2 U3398 ( .A1(n25914), .A2(n28231), .B1(n26254), .B2(n24888), .ZN(
        n22601) );
  OAI22_X2 U3400 ( .A1(n25935), .A2(n28232), .B1(n26254), .B2(n24889), .ZN(
        n22602) );
  OAI22_X2 U3402 ( .A1(n25947), .A2(n28233), .B1(n26254), .B2(n24844), .ZN(
        n22603) );
  OAI22_X2 U3404 ( .A1(n25917), .A2(n28234), .B1(n26254), .B2(n25916), .ZN(
        n22604) );
  OAI22_X2 U3406 ( .A1(n25938), .A2(n28235), .B1(n26254), .B2(n24841), .ZN(
        n22605) );
  OAI22_X2 U3408 ( .A1(n25950), .A2(n28236), .B1(n26254), .B2(n25949), .ZN(
        n22606) );
  OAI22_X2 U3410 ( .A1(n25955), .A2(n26254), .B1(n25957), .B2(n28237), .ZN(
        n22607) );
  OAI22_X2 U3413 ( .A1(n25926), .A2(n28222), .B1(n26255), .B2(n24838), .ZN(
        n22608) );
  OAI22_X2 U3415 ( .A1(n25914), .A2(n28223), .B1(n26255), .B2(n24888), .ZN(
        n22609) );
  OAI22_X2 U3417 ( .A1(n25935), .A2(n28224), .B1(n26255), .B2(n24889), .ZN(
        n22610) );
  OAI22_X2 U3419 ( .A1(n25947), .A2(n28225), .B1(n26255), .B2(n24844), .ZN(
        n22611) );
  OAI22_X2 U3421 ( .A1(n25917), .A2(n28226), .B1(n26255), .B2(n25916), .ZN(
        n22612) );
  OAI22_X2 U3423 ( .A1(n25938), .A2(n28227), .B1(n26255), .B2(n24841), .ZN(
        n22613) );
  OAI22_X2 U3425 ( .A1(n25950), .A2(n28228), .B1(n26255), .B2(n25949), .ZN(
        n22614) );
  OAI22_X2 U3427 ( .A1(n25955), .A2(n26255), .B1(n25956), .B2(n28229), .ZN(
        n22615) );
  OAI22_X2 U3430 ( .A1(n25926), .A2(n28214), .B1(n26256), .B2(n24838), .ZN(
        n22616) );
  OAI22_X2 U3432 ( .A1(n25914), .A2(n28215), .B1(n26256), .B2(n24888), .ZN(
        n22617) );
  OAI22_X2 U3434 ( .A1(n25935), .A2(n28216), .B1(n26256), .B2(n24889), .ZN(
        n22618) );
  OAI22_X2 U3436 ( .A1(n25947), .A2(n28217), .B1(n26256), .B2(n24844), .ZN(
        n22619) );
  OAI22_X2 U3438 ( .A1(n25917), .A2(n28218), .B1(n26256), .B2(n25916), .ZN(
        n22620) );
  OAI22_X2 U3440 ( .A1(n25938), .A2(n28219), .B1(n26256), .B2(n24841), .ZN(
        n22621) );
  OAI22_X2 U3444 ( .A1(n25955), .A2(n26256), .B1(n25956), .B2(n28221), .ZN(
        n22623) );
  OAI22_X2 U3447 ( .A1(n25926), .A2(n28206), .B1(n26257), .B2(n24838), .ZN(
        n22624) );
  OAI22_X2 U3449 ( .A1(n25914), .A2(n28207), .B1(n26257), .B2(n24888), .ZN(
        n22625) );
  OAI22_X2 U3451 ( .A1(n25935), .A2(n28208), .B1(n26257), .B2(n24889), .ZN(
        n22626) );
  OAI22_X2 U3453 ( .A1(n25947), .A2(n28209), .B1(n26257), .B2(n24844), .ZN(
        n22627) );
  OAI22_X2 U3455 ( .A1(n25917), .A2(n28210), .B1(n26257), .B2(n25916), .ZN(
        n22628) );
  OAI22_X2 U3457 ( .A1(n25938), .A2(n28211), .B1(n26257), .B2(n24841), .ZN(
        n22629) );
  OAI22_X2 U3459 ( .A1(n25950), .A2(n28212), .B1(n26257), .B2(n25949), .ZN(
        n22630) );
  OAI22_X2 U3461 ( .A1(n25955), .A2(n26257), .B1(n25957), .B2(n28213), .ZN(
        n22631) );
  OAI22_X2 U3464 ( .A1(n25927), .A2(n28198), .B1(n26258), .B2(n25925), .ZN(
        n22632) );
  OAI22_X2 U3466 ( .A1(n25915), .A2(n28199), .B1(n26258), .B2(n25913), .ZN(
        n22633) );
  OAI22_X2 U3468 ( .A1(n25936), .A2(n28200), .B1(n26258), .B2(n25934), .ZN(
        n22634) );
  OAI22_X2 U3470 ( .A1(n25948), .A2(n28201), .B1(n26258), .B2(n25946), .ZN(
        n22635) );
  OAI22_X2 U3472 ( .A1(n25918), .A2(n28202), .B1(n26258), .B2(n25916), .ZN(
        n22636) );
  OAI22_X2 U3474 ( .A1(n25939), .A2(n28203), .B1(n26258), .B2(n25937), .ZN(
        n22637) );
  OAI22_X2 U3476 ( .A1(n25951), .A2(n28204), .B1(n26258), .B2(n25949), .ZN(
        n22638) );
  OAI22_X2 U3481 ( .A1(n25927), .A2(n28190), .B1(n26259), .B2(n25925), .ZN(
        n22640) );
  OAI22_X2 U3483 ( .A1(n25915), .A2(n28191), .B1(n26259), .B2(n25913), .ZN(
        n22641) );
  OAI22_X2 U3485 ( .A1(n25936), .A2(n28192), .B1(n26259), .B2(n25934), .ZN(
        n22642) );
  OAI22_X2 U3487 ( .A1(n25948), .A2(n28193), .B1(n26259), .B2(n25946), .ZN(
        n22643) );
  OAI22_X2 U3489 ( .A1(n25918), .A2(n28194), .B1(n26259), .B2(n25916), .ZN(
        n22644) );
  OAI22_X2 U3491 ( .A1(n25939), .A2(n28195), .B1(n26259), .B2(n25937), .ZN(
        n22645) );
  OAI22_X2 U3493 ( .A1(n25951), .A2(n28196), .B1(n26259), .B2(n25949), .ZN(
        n22646) );
  OAI22_X2 U3495 ( .A1(n25955), .A2(n26259), .B1(n25957), .B2(n28197), .ZN(
        n22647) );
  OAI22_X2 U3498 ( .A1(n25927), .A2(n28182), .B1(n26260), .B2(n25925), .ZN(
        n22648) );
  OAI22_X2 U3500 ( .A1(n25915), .A2(n28183), .B1(n26260), .B2(n25913), .ZN(
        n22649) );
  OAI22_X2 U3502 ( .A1(n25936), .A2(n28184), .B1(n26260), .B2(n25934), .ZN(
        n22650) );
  OAI22_X2 U3504 ( .A1(n25948), .A2(n28185), .B1(n26260), .B2(n25946), .ZN(
        n22651) );
  OAI22_X2 U3506 ( .A1(n25918), .A2(n28186), .B1(n26260), .B2(n24834), .ZN(
        n22652) );
  OAI22_X2 U3508 ( .A1(n25939), .A2(n28187), .B1(n26260), .B2(n25937), .ZN(
        n22653) );
  OAI22_X2 U3510 ( .A1(n25951), .A2(n28188), .B1(n26260), .B2(n25949), .ZN(
        n22654) );
  OAI22_X2 U3515 ( .A1(n25927), .A2(n28174), .B1(n26261), .B2(n25925), .ZN(
        n22656) );
  OAI22_X2 U3517 ( .A1(n25915), .A2(n28175), .B1(n26261), .B2(n25913), .ZN(
        n22657) );
  OAI22_X2 U3519 ( .A1(n25936), .A2(n28176), .B1(n26261), .B2(n25934), .ZN(
        n22658) );
  OAI22_X2 U3521 ( .A1(n25948), .A2(n28177), .B1(n26261), .B2(n25946), .ZN(
        n22659) );
  OAI22_X2 U3523 ( .A1(n25918), .A2(n28178), .B1(n26261), .B2(n25916), .ZN(
        n22660) );
  OAI22_X2 U3525 ( .A1(n25939), .A2(n28179), .B1(n26261), .B2(n25937), .ZN(
        n22661) );
  OAI22_X2 U3527 ( .A1(n25951), .A2(n28180), .B1(n26261), .B2(n25949), .ZN(
        n22662) );
  OAI22_X2 U3529 ( .A1(n25955), .A2(n26261), .B1(n25957), .B2(n28181), .ZN(
        n22663) );
  OAI22_X2 U3532 ( .A1(n25927), .A2(n28166), .B1(n26262), .B2(n25925), .ZN(
        n22664) );
  OAI22_X2 U3534 ( .A1(n25915), .A2(n28167), .B1(n26262), .B2(n25913), .ZN(
        n22665) );
  OAI22_X2 U3536 ( .A1(n25936), .A2(n28168), .B1(n26262), .B2(n25934), .ZN(
        n22666) );
  OAI22_X2 U3538 ( .A1(n25948), .A2(n28169), .B1(n26262), .B2(n25946), .ZN(
        n22667) );
  OAI22_X2 U3540 ( .A1(n25918), .A2(n28170), .B1(n26262), .B2(n25916), .ZN(
        n22668) );
  OAI22_X2 U3542 ( .A1(n25939), .A2(n28171), .B1(n26262), .B2(n25937), .ZN(
        n22669) );
  OAI22_X2 U3544 ( .A1(n25951), .A2(n28172), .B1(n26262), .B2(n25949), .ZN(
        n22670) );
  OAI22_X2 U3549 ( .A1(n25927), .A2(n28158), .B1(n26263), .B2(n25925), .ZN(
        n22672) );
  OAI22_X2 U3551 ( .A1(n25915), .A2(n28159), .B1(n26263), .B2(n25913), .ZN(
        n22673) );
  OAI22_X2 U3553 ( .A1(n25936), .A2(n28160), .B1(n26263), .B2(n25934), .ZN(
        n22674) );
  OAI22_X2 U3555 ( .A1(n25948), .A2(n28161), .B1(n26263), .B2(n25946), .ZN(
        n22675) );
  OAI22_X2 U3557 ( .A1(n25918), .A2(n28162), .B1(n26263), .B2(n25916), .ZN(
        n22676) );
  OAI22_X2 U3559 ( .A1(n25939), .A2(n28163), .B1(n26263), .B2(n25937), .ZN(
        n22677) );
  OAI22_X2 U3561 ( .A1(n25951), .A2(n28164), .B1(n26263), .B2(n25949), .ZN(
        n22678) );
  OAI22_X2 U3563 ( .A1(n24846), .A2(n26263), .B1(n25957), .B2(n28165), .ZN(
        n22679) );
  OAI22_X2 U3566 ( .A1(n25927), .A2(n28150), .B1(n26264), .B2(n25925), .ZN(
        n22680) );
  OAI22_X2 U3568 ( .A1(n25915), .A2(n28151), .B1(n26264), .B2(n25913), .ZN(
        n22681) );
  OAI22_X2 U3570 ( .A1(n25936), .A2(n28152), .B1(n26264), .B2(n25934), .ZN(
        n22682) );
  OAI22_X2 U3572 ( .A1(n25948), .A2(n28153), .B1(n26264), .B2(n25946), .ZN(
        n22683) );
  OAI22_X2 U3574 ( .A1(n25918), .A2(n28154), .B1(n26264), .B2(n24834), .ZN(
        n22684) );
  OAI22_X2 U3576 ( .A1(n25939), .A2(n28155), .B1(n26264), .B2(n25937), .ZN(
        n22685) );
  OAI22_X2 U3578 ( .A1(n25951), .A2(n28156), .B1(n26264), .B2(n25949), .ZN(
        n22686) );
  OAI22_X2 U3580 ( .A1(n24846), .A2(n26264), .B1(n25957), .B2(n28157), .ZN(
        n22687) );
  OAI22_X2 U3583 ( .A1(n25927), .A2(n28142), .B1(n26265), .B2(n25925), .ZN(
        n22688) );
  OAI22_X2 U3585 ( .A1(n25915), .A2(n28143), .B1(n26265), .B2(n25913), .ZN(
        n22689) );
  OAI22_X2 U3587 ( .A1(n25936), .A2(n28144), .B1(n26265), .B2(n25934), .ZN(
        n22690) );
  OAI22_X2 U3589 ( .A1(n25948), .A2(n28145), .B1(n26265), .B2(n25946), .ZN(
        n22691) );
  OAI22_X2 U3591 ( .A1(n25918), .A2(n28146), .B1(n26265), .B2(n24834), .ZN(
        n22692) );
  OAI22_X2 U3593 ( .A1(n25939), .A2(n28147), .B1(n26265), .B2(n25937), .ZN(
        n22693) );
  OAI22_X2 U3595 ( .A1(n25951), .A2(n28148), .B1(n26265), .B2(n25949), .ZN(
        n22694) );
  OAI22_X2 U3597 ( .A1(n24846), .A2(n26265), .B1(n25957), .B2(n28149), .ZN(
        n22695) );
  OAI22_X2 U3600 ( .A1(n25927), .A2(n28134), .B1(n26266), .B2(n25925), .ZN(
        n22696) );
  OAI22_X2 U3602 ( .A1(n25915), .A2(n28135), .B1(n26266), .B2(n25913), .ZN(
        n22697) );
  OAI22_X2 U3604 ( .A1(n25936), .A2(n28136), .B1(n26266), .B2(n25934), .ZN(
        n22698) );
  OAI22_X2 U3606 ( .A1(n25948), .A2(n28137), .B1(n26266), .B2(n25946), .ZN(
        n22699) );
  OAI22_X2 U3608 ( .A1(n25918), .A2(n28138), .B1(n26266), .B2(n24834), .ZN(
        n22700) );
  OAI22_X2 U3610 ( .A1(n25939), .A2(n28139), .B1(n26266), .B2(n25937), .ZN(
        n22701) );
  OAI22_X2 U3612 ( .A1(n25951), .A2(n28140), .B1(n26266), .B2(n25949), .ZN(
        n22702) );
  OAI22_X2 U3614 ( .A1(n24846), .A2(n26266), .B1(n25957), .B2(n28141), .ZN(
        n22703) );
  OAI22_X2 U3665 ( .A1(n25953), .A2(n28369), .B1(n26193), .B2(n25952), .ZN(
        n22727) );
  OAI22_X2 U3668 ( .A1(n25923), .A2(n28354), .B1(n26194), .B2(n24837), .ZN(
        n22728) );
  OAI22_X2 U3670 ( .A1(n25911), .A2(n28355), .B1(n26194), .B2(n24835), .ZN(
        n22729) );
  OAI22_X2 U3672 ( .A1(n25932), .A2(n28356), .B1(n26194), .B2(n24840), .ZN(
        n22730) );
  OAI22_X2 U3674 ( .A1(n25944), .A2(n28357), .B1(n26194), .B2(n24843), .ZN(
        n22731) );
  OAI22_X2 U3676 ( .A1(n25920), .A2(n28358), .B1(n26194), .B2(n24836), .ZN(
        n22732) );
  OAI22_X2 U3678 ( .A1(n25941), .A2(n28359), .B1(n26194), .B2(n24842), .ZN(
        n22733) );
  OAI22_X2 U3680 ( .A1(n25929), .A2(n28360), .B1(n26194), .B2(n24839), .ZN(
        n22734) );
  OAI22_X2 U3682 ( .A1(n25953), .A2(n28361), .B1(n26194), .B2(n25952), .ZN(
        n22735) );
  OAI22_X2 U3685 ( .A1(n25923), .A2(n28346), .B1(n26195), .B2(n24837), .ZN(
        n22736) );
  OAI22_X2 U3687 ( .A1(n25911), .A2(n28347), .B1(n26195), .B2(n24835), .ZN(
        n22737) );
  OAI22_X2 U3689 ( .A1(n25932), .A2(n28348), .B1(n26195), .B2(n24840), .ZN(
        n22738) );
  OAI22_X2 U3691 ( .A1(n25944), .A2(n28349), .B1(n26195), .B2(n24843), .ZN(
        n22739) );
  OAI22_X2 U3693 ( .A1(n25920), .A2(n28350), .B1(n26195), .B2(n24836), .ZN(
        n22740) );
  OAI22_X2 U3695 ( .A1(n25941), .A2(n28351), .B1(n26195), .B2(n24842), .ZN(
        n22741) );
  OAI22_X2 U3697 ( .A1(n25929), .A2(n28352), .B1(n26195), .B2(n24839), .ZN(
        n22742) );
  OAI22_X2 U3702 ( .A1(n25923), .A2(n28338), .B1(n26196), .B2(n24837), .ZN(
        n22744) );
  OAI22_X2 U3704 ( .A1(n25911), .A2(n28339), .B1(n26196), .B2(n24835), .ZN(
        n22745) );
  OAI22_X2 U3706 ( .A1(n25932), .A2(n28340), .B1(n26196), .B2(n24840), .ZN(
        n22746) );
  OAI22_X2 U3708 ( .A1(n25944), .A2(n28341), .B1(n26196), .B2(n24843), .ZN(
        n22747) );
  OAI22_X2 U3710 ( .A1(n25920), .A2(n28342), .B1(n26196), .B2(n24836), .ZN(
        n22748) );
  OAI22_X2 U3712 ( .A1(n25941), .A2(n28343), .B1(n26196), .B2(n24842), .ZN(
        n22749) );
  OAI22_X2 U3714 ( .A1(n25929), .A2(n28344), .B1(n26196), .B2(n24839), .ZN(
        n22750) );
  OAI22_X2 U3716 ( .A1(n25953), .A2(n28345), .B1(n26196), .B2(n25952), .ZN(
        n22751) );
  OAI22_X2 U3719 ( .A1(n25923), .A2(n28330), .B1(n26197), .B2(n24837), .ZN(
        n22752) );
  OAI22_X2 U3721 ( .A1(n25911), .A2(n28331), .B1(n26197), .B2(n24835), .ZN(
        n22753) );
  OAI22_X2 U3723 ( .A1(n25932), .A2(n28332), .B1(n26197), .B2(n24840), .ZN(
        n22754) );
  OAI22_X2 U3725 ( .A1(n25944), .A2(n28333), .B1(n26197), .B2(n24843), .ZN(
        n22755) );
  OAI22_X2 U3727 ( .A1(n25920), .A2(n28334), .B1(n26197), .B2(n24836), .ZN(
        n22756) );
  OAI22_X2 U3729 ( .A1(n25941), .A2(n28335), .B1(n26197), .B2(n24842), .ZN(
        n22757) );
  OAI22_X2 U3731 ( .A1(n25929), .A2(n28336), .B1(n26197), .B2(n24839), .ZN(
        n22758) );
  OAI22_X2 U3733 ( .A1(n25953), .A2(n28337), .B1(n26197), .B2(n25952), .ZN(
        n22759) );
  OAI22_X2 U3736 ( .A1(n25924), .A2(n28322), .B1(n26198), .B2(n25922), .ZN(
        n22760) );
  OAI22_X2 U3738 ( .A1(n25912), .A2(n28323), .B1(n26198), .B2(n25910), .ZN(
        n22761) );
  OAI22_X2 U3740 ( .A1(n25933), .A2(n28324), .B1(n26198), .B2(n25931), .ZN(
        n22762) );
  OAI22_X2 U3742 ( .A1(n25945), .A2(n28325), .B1(n26198), .B2(n25943), .ZN(
        n22763) );
  OAI22_X2 U3744 ( .A1(n25921), .A2(n28326), .B1(n26198), .B2(n25919), .ZN(
        n22764) );
  OAI22_X2 U3746 ( .A1(n25942), .A2(n28327), .B1(n26198), .B2(n25940), .ZN(
        n22765) );
  OAI22_X2 U3748 ( .A1(n25930), .A2(n28328), .B1(n26198), .B2(n25928), .ZN(
        n22766) );
  OAI22_X2 U3750 ( .A1(n25954), .A2(n28329), .B1(n26198), .B2(n24864), .ZN(
        n22767) );
  OAI22_X2 U3753 ( .A1(n25924), .A2(n28314), .B1(n26199), .B2(n25922), .ZN(
        n22768) );
  OAI22_X2 U3755 ( .A1(n25912), .A2(n28315), .B1(n26199), .B2(n25910), .ZN(
        n22769) );
  OAI22_X2 U3757 ( .A1(n25933), .A2(n28316), .B1(n26199), .B2(n25931), .ZN(
        n22770) );
  OAI22_X2 U3759 ( .A1(n25945), .A2(n28317), .B1(n26199), .B2(n25943), .ZN(
        n22771) );
  OAI22_X2 U3761 ( .A1(n25921), .A2(n28318), .B1(n26199), .B2(n25919), .ZN(
        n22772) );
  OAI22_X2 U3763 ( .A1(n25942), .A2(n28319), .B1(n26199), .B2(n25940), .ZN(
        n22773) );
  OAI22_X2 U3765 ( .A1(n25930), .A2(n28320), .B1(n26199), .B2(n25928), .ZN(
        n22774) );
  OAI22_X2 U3767 ( .A1(n25954), .A2(n28321), .B1(n26199), .B2(n25952), .ZN(
        n22775) );
  OAI22_X2 U3770 ( .A1(n25924), .A2(n28306), .B1(n26200), .B2(n25922), .ZN(
        n22776) );
  OAI22_X2 U3772 ( .A1(n25912), .A2(n28307), .B1(n26200), .B2(n25910), .ZN(
        n22777) );
  OAI22_X2 U3774 ( .A1(n25933), .A2(n28308), .B1(n26200), .B2(n25931), .ZN(
        n22778) );
  OAI22_X2 U3776 ( .A1(n25945), .A2(n28309), .B1(n26200), .B2(n25943), .ZN(
        n22779) );
  OAI22_X2 U3778 ( .A1(n25921), .A2(n28310), .B1(n26200), .B2(n25919), .ZN(
        n22780) );
  OAI22_X2 U3780 ( .A1(n25942), .A2(n28311), .B1(n26200), .B2(n25940), .ZN(
        n22781) );
  OAI22_X2 U3782 ( .A1(n25930), .A2(n28312), .B1(n26200), .B2(n25928), .ZN(
        n22782) );
  OAI22_X2 U3784 ( .A1(n25954), .A2(n28313), .B1(n26200), .B2(n25952), .ZN(
        n22783) );
  OAI22_X2 U3787 ( .A1(n25924), .A2(n28298), .B1(n26201), .B2(n25922), .ZN(
        n22784) );
  OAI22_X2 U3789 ( .A1(n25912), .A2(n28299), .B1(n26201), .B2(n25910), .ZN(
        n22785) );
  OAI22_X2 U3791 ( .A1(n25933), .A2(n28300), .B1(n26201), .B2(n25931), .ZN(
        n22786) );
  OAI22_X2 U3793 ( .A1(n25945), .A2(n28301), .B1(n26201), .B2(n25943), .ZN(
        n22787) );
  OAI22_X2 U3795 ( .A1(n25921), .A2(n28302), .B1(n26201), .B2(n25919), .ZN(
        n22788) );
  OAI22_X2 U3797 ( .A1(n25942), .A2(n28303), .B1(n26201), .B2(n25940), .ZN(
        n22789) );
  OAI22_X2 U3799 ( .A1(n25930), .A2(n28304), .B1(n26201), .B2(n25928), .ZN(
        n22790) );
  OAI22_X2 U3801 ( .A1(n25954), .A2(n28305), .B1(n26201), .B2(n24864), .ZN(
        n22791) );
  OAI22_X2 U3804 ( .A1(n25924), .A2(n28290), .B1(n26202), .B2(n25922), .ZN(
        n22792) );
  OAI22_X2 U3806 ( .A1(n25912), .A2(n28291), .B1(n26202), .B2(n25910), .ZN(
        n22793) );
  OAI22_X2 U3808 ( .A1(n25933), .A2(n28292), .B1(n26202), .B2(n25931), .ZN(
        n22794) );
  OAI22_X2 U3810 ( .A1(n25945), .A2(n28293), .B1(n26202), .B2(n25943), .ZN(
        n22795) );
  OAI22_X2 U3812 ( .A1(n25921), .A2(n28294), .B1(n26202), .B2(n25919), .ZN(
        n22796) );
  OAI22_X2 U3814 ( .A1(n25942), .A2(n28295), .B1(n26202), .B2(n25940), .ZN(
        n22797) );
  OAI22_X2 U3816 ( .A1(n25930), .A2(n28296), .B1(n26202), .B2(n25928), .ZN(
        n22798) );
  OAI22_X2 U3818 ( .A1(n25954), .A2(n28297), .B1(n26202), .B2(n25952), .ZN(
        n22799) );
  OAI22_X2 U3821 ( .A1(n25924), .A2(n28282), .B1(n26203), .B2(n25922), .ZN(
        n22800) );
  OAI22_X2 U3823 ( .A1(n25912), .A2(n28283), .B1(n26203), .B2(n25910), .ZN(
        n22801) );
  OAI22_X2 U3825 ( .A1(n25933), .A2(n28284), .B1(n26203), .B2(n25931), .ZN(
        n22802) );
  OAI22_X2 U3827 ( .A1(n25945), .A2(n28285), .B1(n26203), .B2(n25943), .ZN(
        n22803) );
  OAI22_X2 U3829 ( .A1(n25921), .A2(n28286), .B1(n26203), .B2(n25919), .ZN(
        n22804) );
  OAI22_X2 U3831 ( .A1(n25942), .A2(n28287), .B1(n26203), .B2(n25940), .ZN(
        n22805) );
  OAI22_X2 U3833 ( .A1(n25930), .A2(n28288), .B1(n26203), .B2(n25928), .ZN(
        n22806) );
  OAI22_X2 U3835 ( .A1(n25954), .A2(n28289), .B1(n26203), .B2(n24864), .ZN(
        n22807) );
  OAI22_X2 U3838 ( .A1(n25924), .A2(n28274), .B1(n26204), .B2(n25922), .ZN(
        n22808) );
  OAI22_X2 U3840 ( .A1(n25912), .A2(n28275), .B1(n26204), .B2(n25910), .ZN(
        n22809) );
  OAI22_X2 U3842 ( .A1(n25933), .A2(n28276), .B1(n26204), .B2(n25931), .ZN(
        n22810) );
  OAI22_X2 U3844 ( .A1(n25945), .A2(n28277), .B1(n26204), .B2(n25943), .ZN(
        n22811) );
  OAI22_X2 U3846 ( .A1(n25921), .A2(n28278), .B1(n26204), .B2(n25919), .ZN(
        n22812) );
  OAI22_X2 U3848 ( .A1(n25942), .A2(n28279), .B1(n26204), .B2(n25940), .ZN(
        n22813) );
  OAI22_X2 U3850 ( .A1(n25930), .A2(n28280), .B1(n26204), .B2(n25928), .ZN(
        n22814) );
  OAI22_X2 U3852 ( .A1(n25954), .A2(n28281), .B1(n26204), .B2(n24864), .ZN(
        n22815) );
  OAI22_X2 U3855 ( .A1(n25924), .A2(n28266), .B1(n26205), .B2(n25922), .ZN(
        n22816) );
  OAI22_X2 U3857 ( .A1(n25912), .A2(n28267), .B1(n26205), .B2(n25910), .ZN(
        n22817) );
  OAI22_X2 U3859 ( .A1(n25933), .A2(n28268), .B1(n26205), .B2(n25931), .ZN(
        n22818) );
  OAI22_X2 U3861 ( .A1(n25945), .A2(n28269), .B1(n26205), .B2(n25943), .ZN(
        n22819) );
  OAI22_X2 U3863 ( .A1(n25921), .A2(n28270), .B1(n26205), .B2(n25919), .ZN(
        n22820) );
  OAI22_X2 U3865 ( .A1(n25942), .A2(n28271), .B1(n26205), .B2(n25940), .ZN(
        n22821) );
  OAI22_X2 U3867 ( .A1(n25930), .A2(n28272), .B1(n26205), .B2(n25928), .ZN(
        n22822) );
  OAI22_X2 U3869 ( .A1(n25954), .A2(n28273), .B1(n26205), .B2(n24864), .ZN(
        n22823) );
  OAI22_X2 U3872 ( .A1(n25924), .A2(n28258), .B1(n26206), .B2(n25922), .ZN(
        n22824) );
  OAI22_X2 U3874 ( .A1(n25912), .A2(n28259), .B1(n26206), .B2(n25910), .ZN(
        n22825) );
  OAI22_X2 U3876 ( .A1(n25933), .A2(n28260), .B1(n26206), .B2(n25931), .ZN(
        n22826) );
  OAI22_X2 U3878 ( .A1(n25945), .A2(n28261), .B1(n26206), .B2(n25943), .ZN(
        n22827) );
  OAI22_X2 U3880 ( .A1(n25921), .A2(n28262), .B1(n26206), .B2(n25919), .ZN(
        n22828) );
  OAI22_X2 U3882 ( .A1(n25942), .A2(n28263), .B1(n26206), .B2(n25940), .ZN(
        n22829) );
  OAI22_X2 U3884 ( .A1(n25930), .A2(n28264), .B1(n26206), .B2(n25928), .ZN(
        n22830) );
  OAI22_X2 U3886 ( .A1(n25954), .A2(n28265), .B1(n26206), .B2(n24864), .ZN(
        n22831) );
  OAI22_X2 U3902 ( .A1(n25927), .A2(n28501), .B1(n26207), .B2(n25925), .ZN(
        n22838) );
  OAI22_X2 U3904 ( .A1(n25915), .A2(n28502), .B1(n26207), .B2(n25913), .ZN(
        n22839) );
  OAI22_X2 U3906 ( .A1(n25936), .A2(n28503), .B1(n26207), .B2(n25934), .ZN(
        n22840) );
  OAI22_X2 U3908 ( .A1(n25948), .A2(n28504), .B1(n26207), .B2(n25946), .ZN(
        n22841) );
  OAI22_X2 U3910 ( .A1(n25939), .A2(n28505), .B1(n26207), .B2(n25937), .ZN(
        n22842) );
  OAI22_X2 U3912 ( .A1(n25951), .A2(n28506), .B1(n26207), .B2(n25949), .ZN(
        n22843) );
  OAI22_X2 U3915 ( .A1(n25927), .A2(n28494), .B1(n26208), .B2(n25925), .ZN(
        n22844) );
  OAI22_X2 U3917 ( .A1(n25915), .A2(n28495), .B1(n26208), .B2(n25913), .ZN(
        n22845) );
  OAI22_X2 U3919 ( .A1(n25936), .A2(n28496), .B1(n26208), .B2(n25934), .ZN(
        n22846) );
  OAI22_X2 U3921 ( .A1(n25948), .A2(n28497), .B1(n26208), .B2(n25946), .ZN(
        n22847) );
  OAI22_X2 U3923 ( .A1(n25939), .A2(n28498), .B1(n26208), .B2(n25937), .ZN(
        n22848) );
  OAI22_X2 U3925 ( .A1(n25951), .A2(n28499), .B1(n26208), .B2(n25949), .ZN(
        n22849) );
  OAI22_X2 U3928 ( .A1(n25927), .A2(n28487), .B1(n26209), .B2(n25925), .ZN(
        n22850) );
  OAI22_X2 U3930 ( .A1(n25915), .A2(n28488), .B1(n26209), .B2(n25913), .ZN(
        n22851) );
  OAI22_X2 U3932 ( .A1(n25936), .A2(n28489), .B1(n26209), .B2(n25934), .ZN(
        n22852) );
  OAI22_X2 U3934 ( .A1(n25948), .A2(n28490), .B1(n26209), .B2(n25946), .ZN(
        n22853) );
  OAI22_X2 U3936 ( .A1(n25939), .A2(n28491), .B1(n26209), .B2(n25937), .ZN(
        n22854) );
  OAI22_X2 U3938 ( .A1(n25951), .A2(n28492), .B1(n26209), .B2(n25949), .ZN(
        n22855) );
  OAI22_X2 U3941 ( .A1(n25927), .A2(n28480), .B1(n26210), .B2(n25925), .ZN(
        n22856) );
  OAI22_X2 U3943 ( .A1(n25915), .A2(n28481), .B1(n26210), .B2(n25913), .ZN(
        n22857) );
  OAI22_X2 U3945 ( .A1(n25936), .A2(n28482), .B1(n26210), .B2(n25934), .ZN(
        n22858) );
  OAI22_X2 U3947 ( .A1(n25948), .A2(n28483), .B1(n26210), .B2(n25946), .ZN(
        n22859) );
  OAI22_X2 U3949 ( .A1(n25939), .A2(n28484), .B1(n26210), .B2(n25937), .ZN(
        n22860) );
  OAI22_X2 U3954 ( .A1(n25927), .A2(n28473), .B1(n26211), .B2(n25925), .ZN(
        n22862) );
  OAI22_X2 U3956 ( .A1(n25915), .A2(n28474), .B1(n26211), .B2(n25913), .ZN(
        n22863) );
  OAI22_X2 U3958 ( .A1(n25936), .A2(n28475), .B1(n26211), .B2(n25934), .ZN(
        n22864) );
  OAI22_X2 U3960 ( .A1(n25948), .A2(n28476), .B1(n26211), .B2(n25946), .ZN(
        n22865) );
  OAI22_X2 U3962 ( .A1(n25939), .A2(n28477), .B1(n26211), .B2(n25937), .ZN(
        n22866) );
  OAI22_X2 U3967 ( .A1(n25927), .A2(n28466), .B1(n26212), .B2(n25925), .ZN(
        n22868) );
  OAI22_X2 U3969 ( .A1(n25915), .A2(n28467), .B1(n26212), .B2(n25913), .ZN(
        n22869) );
  OAI22_X2 U3971 ( .A1(n25936), .A2(n28468), .B1(n26212), .B2(n25934), .ZN(
        n22870) );
  OAI22_X2 U3973 ( .A1(n25948), .A2(n28469), .B1(n26212), .B2(n25946), .ZN(
        n22871) );
  OAI22_X2 U3975 ( .A1(n25939), .A2(n28470), .B1(n26212), .B2(n25937), .ZN(
        n22872) );
  OAI22_X2 U3977 ( .A1(n25951), .A2(n28471), .B1(n26212), .B2(n24845), .ZN(
        n22873) );
  OAI22_X2 U3980 ( .A1(n25927), .A2(n28459), .B1(n26213), .B2(n25925), .ZN(
        n22874) );
  OAI22_X2 U3982 ( .A1(n25915), .A2(n28460), .B1(n26213), .B2(n25913), .ZN(
        n22875) );
  OAI22_X2 U3984 ( .A1(n25936), .A2(n28461), .B1(n26213), .B2(n25934), .ZN(
        n22876) );
  OAI22_X2 U3986 ( .A1(n25948), .A2(n28462), .B1(n26213), .B2(n25946), .ZN(
        n22877) );
  OAI22_X2 U3988 ( .A1(n25939), .A2(n28463), .B1(n26213), .B2(n25937), .ZN(
        n22878) );
  OAI22_X2 U3990 ( .A1(n25951), .A2(n28464), .B1(n26213), .B2(n24845), .ZN(
        n22879) );
  OAI22_X2 U3993 ( .A1(n25927), .A2(n28452), .B1(n26214), .B2(n25925), .ZN(
        n22880) );
  OAI22_X2 U3995 ( .A1(n25915), .A2(n28453), .B1(n26214), .B2(n25913), .ZN(
        n22881) );
  OAI22_X2 U3997 ( .A1(n25936), .A2(n28454), .B1(n26214), .B2(n25934), .ZN(
        n22882) );
  OAI22_X2 U3999 ( .A1(n25948), .A2(n28455), .B1(n26214), .B2(n25946), .ZN(
        n22883) );
  OAI22_X2 U4001 ( .A1(n25939), .A2(n28456), .B1(n26214), .B2(n25937), .ZN(
        n22884) );
  OAI22_X2 U4003 ( .A1(n25951), .A2(n28457), .B1(n26214), .B2(n24845), .ZN(
        n22885) );
  OAI22_X2 U4006 ( .A1(n25927), .A2(n28445), .B1(n26215), .B2(n25925), .ZN(
        n22886) );
  OAI22_X2 U4008 ( .A1(n25915), .A2(n28446), .B1(n26215), .B2(n25913), .ZN(
        n22887) );
  OAI22_X2 U4010 ( .A1(n25936), .A2(n28447), .B1(n26215), .B2(n25934), .ZN(
        n22888) );
  OAI22_X2 U4012 ( .A1(n25948), .A2(n28448), .B1(n26215), .B2(n25946), .ZN(
        n22889) );
  OAI22_X2 U4014 ( .A1(n25939), .A2(n28449), .B1(n26215), .B2(n25937), .ZN(
        n22890) );
  OAI22_X2 U4016 ( .A1(n25951), .A2(n28450), .B1(n26215), .B2(n24845), .ZN(
        n22891) );
  OAI22_X2 U4019 ( .A1(n25927), .A2(n28438), .B1(n26216), .B2(n25925), .ZN(
        n22892) );
  OAI22_X2 U4021 ( .A1(n25915), .A2(n28439), .B1(n26216), .B2(n25913), .ZN(
        n22893) );
  OAI22_X2 U4023 ( .A1(n25936), .A2(n28440), .B1(n26216), .B2(n25934), .ZN(
        n22894) );
  OAI22_X2 U4025 ( .A1(n25948), .A2(n28441), .B1(n26216), .B2(n25946), .ZN(
        n22895) );
  OAI22_X2 U4027 ( .A1(n25939), .A2(n28442), .B1(n26216), .B2(n25937), .ZN(
        n22896) );
  OAI22_X2 U4029 ( .A1(n25951), .A2(n28443), .B1(n26216), .B2(n24845), .ZN(
        n22897) );
  OAI22_X2 U4032 ( .A1(n25927), .A2(n28431), .B1(n26217), .B2(n25925), .ZN(
        n22898) );
  OAI22_X2 U4034 ( .A1(n25915), .A2(n28432), .B1(n26217), .B2(n25913), .ZN(
        n22899) );
  OAI22_X2 U4036 ( .A1(n25936), .A2(n28433), .B1(n26217), .B2(n25934), .ZN(
        n22900) );
  OAI22_X2 U4038 ( .A1(n25948), .A2(n28434), .B1(n26217), .B2(n25946), .ZN(
        n22901) );
  OAI22_X2 U4040 ( .A1(n25939), .A2(n28435), .B1(n26217), .B2(n25937), .ZN(
        n22902) );
  OAI22_X2 U4042 ( .A1(n25951), .A2(n28436), .B1(n26217), .B2(n24845), .ZN(
        n22903) );
  OAI22_X2 U4045 ( .A1(n25927), .A2(n28419), .B1(n26218), .B2(n25925), .ZN(
        n22904) );
  OAI22_X2 U4047 ( .A1(n25915), .A2(n28420), .B1(n26218), .B2(n25913), .ZN(
        n22905) );
  OAI22_X2 U4049 ( .A1(n25936), .A2(n28421), .B1(n26218), .B2(n25934), .ZN(
        n22906) );
  OAI22_X2 U4051 ( .A1(n25948), .A2(n28422), .B1(n26218), .B2(n25946), .ZN(
        n22907) );
  OAI22_X2 U4053 ( .A1(n25939), .A2(n28423), .B1(n26218), .B2(n25937), .ZN(
        n22908) );
  OAI22_X2 U4055 ( .A1(n25951), .A2(n28424), .B1(n26218), .B2(n24845), .ZN(
        n22909) );
  OAI22_X2 U4058 ( .A1(n25927), .A2(n28407), .B1(n26219), .B2(n25925), .ZN(
        n22910) );
  OAI22_X2 U4060 ( .A1(n25915), .A2(n28408), .B1(n26219), .B2(n25913), .ZN(
        n22911) );
  OAI22_X2 U4062 ( .A1(n25936), .A2(n28409), .B1(n26219), .B2(n25934), .ZN(
        n22912) );
  OAI22_X2 U4064 ( .A1(n25948), .A2(n28410), .B1(n26219), .B2(n25946), .ZN(
        n22913) );
  OAI22_X2 U4066 ( .A1(n25939), .A2(n28411), .B1(n26219), .B2(n25937), .ZN(
        n22914) );
  OAI22_X2 U4068 ( .A1(n25951), .A2(n28412), .B1(n26219), .B2(n24845), .ZN(
        n22915) );
  OAI22_X2 U4071 ( .A1(n25927), .A2(n28395), .B1(n26220), .B2(n25925), .ZN(
        n22916) );
  OAI22_X2 U4073 ( .A1(n25915), .A2(n28396), .B1(n26220), .B2(n25913), .ZN(
        n22917) );
  OAI22_X2 U4075 ( .A1(n25936), .A2(n28397), .B1(n26220), .B2(n25934), .ZN(
        n22918) );
  OAI22_X2 U4077 ( .A1(n25948), .A2(n28398), .B1(n26220), .B2(n25946), .ZN(
        n22919) );
  OAI22_X2 U4079 ( .A1(n25939), .A2(n28399), .B1(n26220), .B2(n25937), .ZN(
        n22920) );
  OAI22_X2 U4081 ( .A1(n25951), .A2(n28400), .B1(n26220), .B2(n24845), .ZN(
        n22921) );
  OAI22_X2 U4084 ( .A1(n25927), .A2(n28383), .B1(n26221), .B2(n25925), .ZN(
        n22922) );
  OAI22_X2 U4088 ( .A1(n25915), .A2(n28384), .B1(n26221), .B2(n25913), .ZN(
        n22923) );
  OAI22_X2 U4092 ( .A1(n25936), .A2(n28385), .B1(n26221), .B2(n25934), .ZN(
        n22924) );
  OAI22_X2 U4096 ( .A1(n25948), .A2(n28386), .B1(n26221), .B2(n25946), .ZN(
        n22925) );
  NOR2_X2 U4100 ( .A1(n24887), .A2(n22403), .ZN(n12056) );
  OAI22_X2 U4101 ( .A1(n25939), .A2(n28387), .B1(n26221), .B2(n25937), .ZN(
        n22926) );
  OAI22_X2 U4105 ( .A1(n25951), .A2(n28388), .B1(n26221), .B2(n24845), .ZN(
        n22927) );
  OAI22_X2 U4131 ( .A1(n25924), .A2(n28681), .B1(n26237), .B2(n25922), .ZN(
        n22938) );
  OAI22_X2 U4133 ( .A1(n25912), .A2(n28682), .B1(n26237), .B2(n25910), .ZN(
        n22939) );
  OAI22_X2 U4135 ( .A1(n25933), .A2(n28683), .B1(n26237), .B2(n25931), .ZN(
        n22940) );
  OAI22_X2 U4137 ( .A1(n25945), .A2(n28684), .B1(n26237), .B2(n25943), .ZN(
        n22941) );
  OAI22_X2 U4139 ( .A1(n25918), .A2(n28685), .B1(n26237), .B2(n24834), .ZN(
        n22942) );
  OAI22_X2 U4141 ( .A1(n25921), .A2(n28686), .B1(n26237), .B2(n25919), .ZN(
        n22943) );
  OAI22_X2 U4143 ( .A1(n25942), .A2(n28687), .B1(n26237), .B2(n25940), .ZN(
        n22944) );
  OAI22_X2 U4145 ( .A1(n25930), .A2(n28688), .B1(n26237), .B2(n25928), .ZN(
        n22945) );
  OAI22_X2 U4147 ( .A1(n25954), .A2(n28689), .B1(n25952), .B2(n26237), .ZN(
        n22946) );
  OAI22_X2 U4149 ( .A1(n24846), .A2(n26237), .B1(n25957), .B2(n28690), .ZN(
        n22947) );
  OAI22_X2 U4152 ( .A1(n25924), .A2(n28670), .B1(n26238), .B2(n25922), .ZN(
        n22948) );
  OAI22_X2 U4154 ( .A1(n25912), .A2(n28671), .B1(n26238), .B2(n25910), .ZN(
        n22949) );
  OAI22_X2 U4156 ( .A1(n25933), .A2(n28672), .B1(n26238), .B2(n25931), .ZN(
        n22950) );
  OAI22_X2 U4158 ( .A1(n25945), .A2(n28673), .B1(n26238), .B2(n25943), .ZN(
        n22951) );
  OAI22_X2 U4160 ( .A1(n25918), .A2(n28674), .B1(n26238), .B2(n24834), .ZN(
        n22952) );
  OAI22_X2 U4162 ( .A1(n25921), .A2(n28675), .B1(n26238), .B2(n25919), .ZN(
        n22953) );
  OAI22_X2 U4164 ( .A1(n25942), .A2(n28676), .B1(n26238), .B2(n25940), .ZN(
        n22954) );
  OAI22_X2 U4166 ( .A1(n25930), .A2(n28677), .B1(n26238), .B2(n25928), .ZN(
        n22955) );
  OAI22_X2 U4168 ( .A1(n25954), .A2(n28678), .B1(n25952), .B2(n26238), .ZN(
        n22956) );
  OAI22_X2 U4170 ( .A1(n24846), .A2(n26238), .B1(n25957), .B2(n28679), .ZN(
        n22957) );
  OAI22_X2 U4173 ( .A1(n25924), .A2(n28659), .B1(n26239), .B2(n25922), .ZN(
        n22958) );
  OAI22_X2 U4175 ( .A1(n25912), .A2(n28660), .B1(n26239), .B2(n25910), .ZN(
        n22959) );
  OAI22_X2 U4177 ( .A1(n25933), .A2(n28661), .B1(n26239), .B2(n25931), .ZN(
        n22960) );
  OAI22_X2 U4179 ( .A1(n25945), .A2(n28662), .B1(n26239), .B2(n25943), .ZN(
        n22961) );
  OAI22_X2 U4181 ( .A1(n25918), .A2(n28663), .B1(n26239), .B2(n24834), .ZN(
        n22962) );
  OAI22_X2 U4183 ( .A1(n25921), .A2(n28664), .B1(n26239), .B2(n25919), .ZN(
        n22963) );
  OAI22_X2 U4185 ( .A1(n25942), .A2(n28665), .B1(n26239), .B2(n25940), .ZN(
        n22964) );
  OAI22_X2 U4187 ( .A1(n25930), .A2(n28666), .B1(n26239), .B2(n25928), .ZN(
        n22965) );
  OAI22_X2 U4189 ( .A1(n25954), .A2(n28667), .B1(n25952), .B2(n26239), .ZN(
        n22966) );
  OAI22_X2 U4191 ( .A1(n24846), .A2(n26239), .B1(n25957), .B2(n28668), .ZN(
        n22967) );
  OAI22_X2 U4194 ( .A1(n25924), .A2(n28648), .B1(n26240), .B2(n25922), .ZN(
        n22968) );
  OAI22_X2 U4196 ( .A1(n25912), .A2(n28649), .B1(n26240), .B2(n25910), .ZN(
        n22969) );
  OAI22_X2 U4198 ( .A1(n25933), .A2(n28650), .B1(n26240), .B2(n25931), .ZN(
        n22970) );
  OAI22_X2 U4200 ( .A1(n25945), .A2(n28651), .B1(n26240), .B2(n25943), .ZN(
        n22971) );
  OAI22_X2 U4202 ( .A1(n25918), .A2(n28652), .B1(n26240), .B2(n25916), .ZN(
        n22972) );
  OAI22_X2 U4204 ( .A1(n25921), .A2(n28653), .B1(n26240), .B2(n25919), .ZN(
        n22973) );
  OAI22_X2 U4206 ( .A1(n25942), .A2(n28654), .B1(n26240), .B2(n25940), .ZN(
        n22974) );
  OAI22_X2 U4208 ( .A1(n25930), .A2(n28655), .B1(n26240), .B2(n25928), .ZN(
        n22975) );
  OAI22_X2 U4210 ( .A1(n25954), .A2(n28656), .B1(n25952), .B2(n26240), .ZN(
        n22976) );
  OAI22_X2 U4212 ( .A1(n25955), .A2(n26240), .B1(n25957), .B2(n28657), .ZN(
        n22977) );
  OAI22_X2 U4215 ( .A1(n25924), .A2(n28637), .B1(n26241), .B2(n25922), .ZN(
        n22978) );
  OAI22_X2 U4217 ( .A1(n25912), .A2(n28638), .B1(n26241), .B2(n25910), .ZN(
        n22979) );
  OAI22_X2 U4219 ( .A1(n25933), .A2(n28639), .B1(n26241), .B2(n25931), .ZN(
        n22980) );
  OAI22_X2 U4221 ( .A1(n25945), .A2(n28640), .B1(n26241), .B2(n25943), .ZN(
        n22981) );
  OAI22_X2 U4223 ( .A1(n25918), .A2(n28641), .B1(n26241), .B2(n25916), .ZN(
        n22982) );
  OAI22_X2 U4225 ( .A1(n25921), .A2(n28642), .B1(n26241), .B2(n25919), .ZN(
        n22983) );
  OAI22_X2 U4227 ( .A1(n25942), .A2(n28643), .B1(n26241), .B2(n25940), .ZN(
        n22984) );
  OAI22_X2 U4229 ( .A1(n25930), .A2(n28644), .B1(n26241), .B2(n25928), .ZN(
        n22985) );
  OAI22_X2 U4231 ( .A1(n25954), .A2(n28645), .B1(n25952), .B2(n26241), .ZN(
        n22986) );
  OAI22_X2 U4233 ( .A1(n25955), .A2(n26241), .B1(n25957), .B2(n28646), .ZN(
        n22987) );
  OAI22_X2 U4236 ( .A1(n25924), .A2(n28626), .B1(n26242), .B2(n25922), .ZN(
        n22988) );
  OAI22_X2 U4238 ( .A1(n25912), .A2(n28627), .B1(n26242), .B2(n25910), .ZN(
        n22989) );
  OAI22_X2 U4240 ( .A1(n25933), .A2(n28628), .B1(n26242), .B2(n25931), .ZN(
        n22990) );
  OAI22_X2 U4242 ( .A1(n25945), .A2(n28629), .B1(n26242), .B2(n25943), .ZN(
        n22991) );
  OAI22_X2 U4244 ( .A1(n25918), .A2(n28630), .B1(n26242), .B2(n25916), .ZN(
        n22992) );
  OAI22_X2 U4246 ( .A1(n25921), .A2(n28631), .B1(n26242), .B2(n25919), .ZN(
        n22993) );
  OAI22_X2 U4248 ( .A1(n25942), .A2(n28632), .B1(n26242), .B2(n25940), .ZN(
        n22994) );
  OAI22_X2 U4250 ( .A1(n25930), .A2(n28633), .B1(n26242), .B2(n25928), .ZN(
        n22995) );
  OAI22_X2 U4252 ( .A1(n25954), .A2(n28634), .B1(n25952), .B2(n26242), .ZN(
        n22996) );
  OAI22_X2 U4254 ( .A1(n25955), .A2(n26242), .B1(n25957), .B2(n28635), .ZN(
        n22997) );
  OAI22_X2 U4257 ( .A1(n25924), .A2(n28615), .B1(n26243), .B2(n25922), .ZN(
        n22998) );
  OAI22_X2 U4259 ( .A1(n25912), .A2(n28616), .B1(n26243), .B2(n25910), .ZN(
        n22999) );
  OAI22_X2 U4261 ( .A1(n25933), .A2(n28617), .B1(n26243), .B2(n25931), .ZN(
        n23000) );
  OAI22_X2 U4263 ( .A1(n25945), .A2(n28618), .B1(n26243), .B2(n25943), .ZN(
        n23001) );
  OAI22_X2 U4265 ( .A1(n25918), .A2(n28619), .B1(n26243), .B2(n25916), .ZN(
        n23002) );
  OAI22_X2 U4267 ( .A1(n25921), .A2(n28620), .B1(n26243), .B2(n25919), .ZN(
        n23003) );
  OAI22_X2 U4269 ( .A1(n25942), .A2(n28621), .B1(n26243), .B2(n25940), .ZN(
        n23004) );
  OAI22_X2 U4271 ( .A1(n25930), .A2(n28622), .B1(n26243), .B2(n25928), .ZN(
        n23005) );
  OAI22_X2 U4273 ( .A1(n25954), .A2(n28623), .B1(n25952), .B2(n26243), .ZN(
        n23006) );
  OAI22_X2 U4275 ( .A1(n25955), .A2(n26243), .B1(n25957), .B2(n28624), .ZN(
        n23007) );
  OAI22_X2 U4278 ( .A1(n25924), .A2(n28604), .B1(n26244), .B2(n25922), .ZN(
        n23008) );
  OAI22_X2 U4280 ( .A1(n25912), .A2(n28605), .B1(n26244), .B2(n25910), .ZN(
        n23009) );
  OAI22_X2 U4282 ( .A1(n25933), .A2(n28606), .B1(n26244), .B2(n25931), .ZN(
        n23010) );
  OAI22_X2 U4284 ( .A1(n25945), .A2(n28607), .B1(n26244), .B2(n25943), .ZN(
        n23011) );
  OAI22_X2 U4286 ( .A1(n25918), .A2(n28608), .B1(n26244), .B2(n25916), .ZN(
        n23012) );
  OAI22_X2 U4288 ( .A1(n25921), .A2(n28609), .B1(n26244), .B2(n25919), .ZN(
        n23013) );
  OAI22_X2 U4290 ( .A1(n25942), .A2(n28610), .B1(n26244), .B2(n25940), .ZN(
        n23014) );
  OAI22_X2 U4292 ( .A1(n25930), .A2(n28611), .B1(n26244), .B2(n25928), .ZN(
        n23015) );
  OAI22_X2 U4294 ( .A1(n25954), .A2(n28612), .B1(n25952), .B2(n26244), .ZN(
        n23016) );
  OAI22_X2 U4296 ( .A1(n25955), .A2(n26244), .B1(n25957), .B2(n28613), .ZN(
        n23017) );
  OAI22_X2 U4299 ( .A1(n25924), .A2(n28593), .B1(n26245), .B2(n25922), .ZN(
        n23018) );
  OAI22_X2 U4301 ( .A1(n25912), .A2(n28594), .B1(n26245), .B2(n25910), .ZN(
        n23019) );
  OAI22_X2 U4303 ( .A1(n25933), .A2(n28595), .B1(n26245), .B2(n25931), .ZN(
        n23020) );
  OAI22_X2 U4305 ( .A1(n25945), .A2(n28596), .B1(n26245), .B2(n25943), .ZN(
        n23021) );
  OAI22_X2 U4307 ( .A1(n25918), .A2(n28597), .B1(n26245), .B2(n25916), .ZN(
        n23022) );
  OAI22_X2 U4309 ( .A1(n25921), .A2(n28598), .B1(n26245), .B2(n25919), .ZN(
        n23023) );
  OAI22_X2 U4311 ( .A1(n25942), .A2(n28599), .B1(n26245), .B2(n25940), .ZN(
        n23024) );
  OAI22_X2 U4313 ( .A1(n25930), .A2(n28600), .B1(n26245), .B2(n25928), .ZN(
        n23025) );
  OAI22_X2 U4315 ( .A1(n25954), .A2(n28601), .B1(n25952), .B2(n26245), .ZN(
        n23026) );
  OAI22_X2 U4317 ( .A1(n25955), .A2(n26245), .B1(n25957), .B2(n28602), .ZN(
        n23027) );
  OAI22_X2 U4320 ( .A1(n25924), .A2(n28582), .B1(n26246), .B2(n25922), .ZN(
        n23028) );
  OAI22_X2 U4322 ( .A1(n25912), .A2(n28583), .B1(n26246), .B2(n25910), .ZN(
        n23029) );
  OAI22_X2 U4324 ( .A1(n25933), .A2(n28584), .B1(n26246), .B2(n25931), .ZN(
        n23030) );
  OAI22_X2 U4326 ( .A1(n25945), .A2(n28585), .B1(n26246), .B2(n25943), .ZN(
        n23031) );
  OAI22_X2 U4328 ( .A1(n25918), .A2(n28586), .B1(n26246), .B2(n25916), .ZN(
        n23032) );
  OAI22_X2 U4330 ( .A1(n25921), .A2(n28587), .B1(n26246), .B2(n25919), .ZN(
        n23033) );
  OAI22_X2 U4332 ( .A1(n25942), .A2(n28588), .B1(n26246), .B2(n25940), .ZN(
        n23034) );
  OAI22_X2 U4334 ( .A1(n25930), .A2(n28589), .B1(n26246), .B2(n25928), .ZN(
        n23035) );
  OAI22_X2 U4336 ( .A1(n25954), .A2(n28590), .B1(n25952), .B2(n26246), .ZN(
        n23036) );
  OAI22_X2 U4338 ( .A1(n25955), .A2(n26246), .B1(n25957), .B2(n28591), .ZN(
        n23037) );
  OAI22_X2 U4341 ( .A1(n25924), .A2(n28571), .B1(n26247), .B2(n25922), .ZN(
        n23038) );
  OAI22_X2 U4343 ( .A1(n25912), .A2(n28572), .B1(n26247), .B2(n25910), .ZN(
        n23039) );
  OAI22_X2 U4345 ( .A1(n25933), .A2(n28573), .B1(n26247), .B2(n25931), .ZN(
        n23040) );
  OAI22_X2 U4347 ( .A1(n25945), .A2(n28574), .B1(n26247), .B2(n25943), .ZN(
        n23041) );
  OAI22_X2 U4349 ( .A1(n25918), .A2(n28575), .B1(n26247), .B2(n25916), .ZN(
        n23042) );
  OAI22_X2 U4351 ( .A1(n25921), .A2(n28576), .B1(n26247), .B2(n25919), .ZN(
        n23043) );
  OAI22_X2 U4353 ( .A1(n25942), .A2(n28577), .B1(n26247), .B2(n25940), .ZN(
        n23044) );
  OAI22_X2 U4355 ( .A1(n25930), .A2(n28578), .B1(n26247), .B2(n25928), .ZN(
        n23045) );
  OAI22_X2 U4357 ( .A1(n25954), .A2(n28579), .B1(n25952), .B2(n26247), .ZN(
        n23046) );
  OAI22_X2 U4359 ( .A1(n25955), .A2(n26247), .B1(n25957), .B2(n28580), .ZN(
        n23047) );
  OAI22_X2 U4362 ( .A1(n25924), .A2(n28556), .B1(n26248), .B2(n25922), .ZN(
        n23048) );
  OAI22_X2 U4364 ( .A1(n25912), .A2(n28557), .B1(n26248), .B2(n25910), .ZN(
        n23049) );
  OAI22_X2 U4366 ( .A1(n25933), .A2(n28558), .B1(n26248), .B2(n25931), .ZN(
        n23050) );
  OAI22_X2 U4368 ( .A1(n25945), .A2(n28559), .B1(n26248), .B2(n25943), .ZN(
        n23051) );
  OAI22_X2 U4370 ( .A1(n25918), .A2(n28560), .B1(n26248), .B2(n25916), .ZN(
        n23052) );
  OAI22_X2 U4372 ( .A1(n25921), .A2(n28561), .B1(n26248), .B2(n25919), .ZN(
        n23053) );
  OAI22_X2 U4374 ( .A1(n25942), .A2(n28562), .B1(n26248), .B2(n25940), .ZN(
        n23054) );
  OAI22_X2 U4376 ( .A1(n25930), .A2(n28563), .B1(n26248), .B2(n25928), .ZN(
        n23055) );
  OAI22_X2 U4378 ( .A1(n25954), .A2(n28564), .B1(n25952), .B2(n26248), .ZN(
        n23056) );
  OAI22_X2 U4380 ( .A1(n25955), .A2(n26248), .B1(n25957), .B2(n28565), .ZN(
        n23057) );
  OAI22_X2 U4383 ( .A1(n25924), .A2(n28541), .B1(n26249), .B2(n25922), .ZN(
        n23058) );
  OAI22_X2 U4385 ( .A1(n25912), .A2(n28542), .B1(n26249), .B2(n25910), .ZN(
        n23059) );
  OAI22_X2 U4387 ( .A1(n25933), .A2(n28543), .B1(n26249), .B2(n25931), .ZN(
        n23060) );
  OAI22_X2 U4389 ( .A1(n25945), .A2(n28544), .B1(n26249), .B2(n25943), .ZN(
        n23061) );
  OAI22_X2 U4391 ( .A1(n25918), .A2(n28545), .B1(n26249), .B2(n25916), .ZN(
        n23062) );
  OAI22_X2 U4393 ( .A1(n25921), .A2(n28546), .B1(n26249), .B2(n25919), .ZN(
        n23063) );
  OAI22_X2 U4395 ( .A1(n25942), .A2(n28547), .B1(n26249), .B2(n25940), .ZN(
        n23064) );
  OAI22_X2 U4397 ( .A1(n25930), .A2(n28548), .B1(n26249), .B2(n25928), .ZN(
        n23065) );
  OAI22_X2 U4399 ( .A1(n25954), .A2(n28549), .B1(n25952), .B2(n26249), .ZN(
        n23066) );
  OAI22_X2 U4401 ( .A1(n25955), .A2(n26249), .B1(n25957), .B2(n28550), .ZN(
        n23067) );
  OAI22_X2 U4404 ( .A1(n25924), .A2(n28526), .B1(n26250), .B2(n25922), .ZN(
        n23068) );
  OAI22_X2 U4406 ( .A1(n25912), .A2(n28527), .B1(n26250), .B2(n25910), .ZN(
        n23069) );
  OAI22_X2 U4408 ( .A1(n25933), .A2(n28528), .B1(n26250), .B2(n25931), .ZN(
        n23070) );
  OAI22_X2 U4410 ( .A1(n25945), .A2(n28529), .B1(n26250), .B2(n25943), .ZN(
        n23071) );
  OAI22_X2 U4412 ( .A1(n25918), .A2(n28530), .B1(n26250), .B2(n25916), .ZN(
        n23072) );
  OAI22_X2 U4414 ( .A1(n25921), .A2(n28531), .B1(n26250), .B2(n25919), .ZN(
        n23073) );
  OAI22_X2 U4416 ( .A1(n25942), .A2(n28532), .B1(n26250), .B2(n25940), .ZN(
        n23074) );
  OAI22_X2 U4418 ( .A1(n25930), .A2(n28533), .B1(n26250), .B2(n25928), .ZN(
        n23075) );
  OAI22_X2 U4420 ( .A1(n25954), .A2(n28534), .B1(n25952), .B2(n26250), .ZN(
        n23076) );
  OAI22_X2 U4422 ( .A1(n25955), .A2(n26250), .B1(n25957), .B2(n28535), .ZN(
        n23077) );
  OAI22_X2 U4425 ( .A1(n25924), .A2(n28511), .B1(n26251), .B2(n25922), .ZN(
        n23078) );
  OAI22_X2 U4429 ( .A1(n25912), .A2(n28512), .B1(n26251), .B2(n25910), .ZN(
        n23079) );
  OAI22_X2 U4433 ( .A1(n25933), .A2(n28513), .B1(n26251), .B2(n25931), .ZN(
        n23080) );
  OAI22_X2 U4437 ( .A1(n25945), .A2(n28514), .B1(n26251), .B2(n25943), .ZN(
        n23081) );
  NOR2_X2 U4441 ( .A1(n25253), .A2(n22402), .ZN(n12140) );
  OAI22_X2 U4442 ( .A1(n25918), .A2(n28515), .B1(n26251), .B2(n25916), .ZN(
        n23082) );
  OAI22_X2 U4446 ( .A1(n25921), .A2(n28516), .B1(n26251), .B2(n25919), .ZN(
        n23083) );
  AND3_X2 U4450 ( .A1(n12146), .A2(n25257), .A3(n22401), .ZN(n12058) );
  OAI22_X2 U4451 ( .A1(n25942), .A2(n28517), .B1(n26251), .B2(n25940), .ZN(
        n23084) );
  AND3_X2 U4455 ( .A1(n12146), .A2(n24896), .A3(n22400), .ZN(n12060) );
  OAI22_X2 U4456 ( .A1(n25930), .A2(n28518), .B1(n26251), .B2(n25928), .ZN(
        n23085) );
  OAI22_X2 U4460 ( .A1(n25954), .A2(n28519), .B1(n25952), .B2(n26251), .ZN(
        n23086) );
  NOR2_X2 U4464 ( .A1(n24887), .A2(n25253), .ZN(n12145) );
  AND3_X2 U4465 ( .A1(n22401), .A2(n12146), .A3(n22400), .ZN(n12062) );
  OAI22_X2 U4466 ( .A1(n25955), .A2(n26251), .B1(n25957), .B2(n28520), .ZN(
        n23087) );
  OAI22_X2 U4469 ( .A1(n25961), .A2(n25907), .B1(n12152), .B2(n12153), .ZN(
        n23088) );
  NOR2_X2 U4470 ( .A1(n12154), .A2(n12155), .ZN(n12152) );
  NAND4_X2 U4471 ( .A1(n12156), .A2(n12157), .A3(n12158), .A4(n12159), .ZN(
        n12155) );
  AOI221_X2 U4472 ( .B1(n12160), .B2(n25731), .C1(n12162), .C2(n25244), .A(
        n12164), .ZN(n12159) );
  AOI221_X2 U4476 ( .B1(n12170), .B2(n25730), .C1(n12172), .C2(n25243), .A(
        n12174), .ZN(n12158) );
  OAI22_X2 U4477 ( .A1(n19340), .A2(n12175), .B1(n19314), .B2(n12176), .ZN(
        n12174) );
  AOI221_X2 U4480 ( .B1(n19321), .B2(n12177), .C1(n19312), .C2(n12178), .A(
        n12179), .ZN(n12157) );
  AOI221_X2 U4482 ( .B1(n19320), .B2(n12185), .C1(n19311), .C2(n12186), .A(
        n12187), .ZN(n12156) );
  OAI22_X2 U4483 ( .A1(n12188), .A2(n27957), .B1(n12190), .B2(n27877), .ZN(
        n12187) );
  NAND4_X2 U4484 ( .A1(n12192), .A2(n12193), .A3(n12194), .A4(n12195), .ZN(
        n12154) );
  AOI221_X2 U4485 ( .B1(n19343), .B2(n12196), .C1(n19342), .C2(n12197), .A(
        n12198), .ZN(n12195) );
  AOI221_X2 U4487 ( .B1(n12203), .B2(n25729), .C1(n12205), .C2(n25242), .A(
        n12207), .ZN(n12194) );
  OAI22_X2 U4488 ( .A1(n12208), .A2(n27909), .B1(n12210), .B2(n27925), .ZN(
        n12207) );
  AOI221_X2 U4491 ( .B1(n19326), .B2(n12212), .C1(n19325), .C2(n12213), .A(
        n12214), .ZN(n12193) );
  AOI221_X2 U4493 ( .B1(n12219), .B2(n25728), .C1(n12221), .C2(n25241), .A(
        n12223), .ZN(n12192) );
  OAI22_X2 U4494 ( .A1(n12224), .A2(n28069), .B1(n12226), .B2(n28085), .ZN(
        n12223) );
  OAI22_X2 U4497 ( .A1(n25963), .A2(n25909), .B1(n12228), .B2(n12153), .ZN(
        n23089) );
  NOR2_X2 U4498 ( .A1(n12229), .A2(n12230), .ZN(n12228) );
  NAND4_X2 U4499 ( .A1(n12231), .A2(n12232), .A3(n12233), .A4(n12234), .ZN(
        n12230) );
  AOI221_X2 U4500 ( .B1(n12160), .B2(n25727), .C1(n12162), .C2(n25240), .A(
        n12237), .ZN(n12234) );
  AOI221_X2 U4504 ( .B1(n12170), .B2(n25726), .C1(n12172), .C2(n25239), .A(
        n12242), .ZN(n12233) );
  OAI22_X2 U4505 ( .A1(n19303), .A2(n12175), .B1(n19277), .B2(n12176), .ZN(
        n12242) );
  AOI221_X2 U4508 ( .B1(n19284), .B2(n12177), .C1(n19275), .C2(n12178), .A(
        n12243), .ZN(n12232) );
  AOI221_X2 U4510 ( .B1(n19283), .B2(n12185), .C1(n19274), .C2(n12186), .A(
        n12246), .ZN(n12231) );
  OAI22_X2 U4511 ( .A1(n12188), .A2(n27956), .B1(n12190), .B2(n27876), .ZN(
        n12246) );
  NAND4_X2 U4512 ( .A1(n12249), .A2(n12250), .A3(n12251), .A4(n12252), .ZN(
        n12229) );
  AOI221_X2 U4513 ( .B1(n19306), .B2(n12196), .C1(n19305), .C2(n12197), .A(
        n12253), .ZN(n12252) );
  AOI221_X2 U4515 ( .B1(n12203), .B2(n25725), .C1(n12205), .C2(n25238), .A(
        n12257), .ZN(n12251) );
  OAI22_X2 U4516 ( .A1(n12208), .A2(n27908), .B1(n12210), .B2(n27924), .ZN(
        n12257) );
  AOI221_X2 U4519 ( .B1(n19289), .B2(n12212), .C1(n19288), .C2(n12213), .A(
        n12260), .ZN(n12250) );
  AOI221_X2 U4521 ( .B1(n12219), .B2(n25724), .C1(n12221), .C2(n25237), .A(
        n12264), .ZN(n12249) );
  OAI22_X2 U4522 ( .A1(n12224), .A2(n28068), .B1(n12226), .B2(n28084), .ZN(
        n12264) );
  OAI22_X2 U4525 ( .A1(n25965), .A2(n25907), .B1(n12267), .B2(n25908), .ZN(
        n23090) );
  NOR2_X2 U4526 ( .A1(n12268), .A2(n12269), .ZN(n12267) );
  NAND4_X2 U4527 ( .A1(n12270), .A2(n12271), .A3(n12272), .A4(n12273), .ZN(
        n12269) );
  AOI221_X2 U4528 ( .B1(n12160), .B2(n25723), .C1(n12162), .C2(n25236), .A(
        n12276), .ZN(n12273) );
  AOI221_X2 U4532 ( .B1(n12170), .B2(n25722), .C1(n12172), .C2(n25235), .A(
        n12281), .ZN(n12272) );
  OAI22_X2 U4533 ( .A1(n19266), .A2(n12175), .B1(n19240), .B2(n12176), .ZN(
        n12281) );
  AOI221_X2 U4536 ( .B1(n19247), .B2(n12177), .C1(n19238), .C2(n12178), .A(
        n12282), .ZN(n12271) );
  AOI221_X2 U4538 ( .B1(n19246), .B2(n12185), .C1(n19237), .C2(n12186), .A(
        n12285), .ZN(n12270) );
  OAI22_X2 U4539 ( .A1(n12188), .A2(n27955), .B1(n12190), .B2(n27875), .ZN(
        n12285) );
  NAND4_X2 U4540 ( .A1(n12288), .A2(n12289), .A3(n12290), .A4(n12291), .ZN(
        n12268) );
  AOI221_X2 U4541 ( .B1(n19269), .B2(n12196), .C1(n19268), .C2(n12197), .A(
        n12292), .ZN(n12291) );
  AOI221_X2 U4543 ( .B1(n12203), .B2(n25721), .C1(n12205), .C2(n25234), .A(
        n12296), .ZN(n12290) );
  OAI22_X2 U4544 ( .A1(n12208), .A2(n27907), .B1(n12210), .B2(n27923), .ZN(
        n12296) );
  AOI221_X2 U4547 ( .B1(n19252), .B2(n12212), .C1(n19251), .C2(n12213), .A(
        n12299), .ZN(n12289) );
  AOI221_X2 U4549 ( .B1(n12219), .B2(n25720), .C1(n12221), .C2(n25233), .A(
        n12303), .ZN(n12288) );
  OAI22_X2 U4550 ( .A1(n12224), .A2(n28067), .B1(n12226), .B2(n28083), .ZN(
        n12303) );
  OAI22_X2 U4553 ( .A1(n25967), .A2(n25909), .B1(n12306), .B2(n25908), .ZN(
        n23091) );
  NOR2_X2 U4554 ( .A1(n12307), .A2(n12308), .ZN(n12306) );
  NAND4_X2 U4555 ( .A1(n12309), .A2(n12310), .A3(n12311), .A4(n12312), .ZN(
        n12308) );
  AOI221_X2 U4556 ( .B1(n12160), .B2(n25719), .C1(n12162), .C2(n25232), .A(
        n12315), .ZN(n12312) );
  AOI221_X2 U4560 ( .B1(n12170), .B2(n25718), .C1(n12172), .C2(n25231), .A(
        n12320), .ZN(n12311) );
  OAI22_X2 U4561 ( .A1(n19229), .A2(n12175), .B1(n19203), .B2(n12176), .ZN(
        n12320) );
  AOI221_X2 U4564 ( .B1(n19210), .B2(n12177), .C1(n19201), .C2(n12178), .A(
        n12321), .ZN(n12310) );
  AOI221_X2 U4566 ( .B1(n19209), .B2(n12185), .C1(n19200), .C2(n12186), .A(
        n12324), .ZN(n12309) );
  OAI22_X2 U4567 ( .A1(n12188), .A2(n27954), .B1(n12190), .B2(n27874), .ZN(
        n12324) );
  NAND4_X2 U4568 ( .A1(n12327), .A2(n12328), .A3(n12329), .A4(n12330), .ZN(
        n12307) );
  AOI221_X2 U4569 ( .B1(n19232), .B2(n12196), .C1(n19231), .C2(n12197), .A(
        n12331), .ZN(n12330) );
  AOI221_X2 U4571 ( .B1(n12203), .B2(n25717), .C1(n12205), .C2(n25230), .A(
        n12335), .ZN(n12329) );
  OAI22_X2 U4572 ( .A1(n12208), .A2(n27906), .B1(n12210), .B2(n27922), .ZN(
        n12335) );
  AOI221_X2 U4575 ( .B1(n19215), .B2(n12212), .C1(n19214), .C2(n12213), .A(
        n12338), .ZN(n12328) );
  AOI221_X2 U4577 ( .B1(n12219), .B2(n25716), .C1(n12221), .C2(n25229), .A(
        n12342), .ZN(n12327) );
  OAI22_X2 U4578 ( .A1(n12224), .A2(n28066), .B1(n12226), .B2(n28082), .ZN(
        n12342) );
  NAND4_X2 U4583 ( .A1(n12348), .A2(n12349), .A3(n12350), .A4(n12351), .ZN(
        n12347) );
  AOI221_X2 U4584 ( .B1(n12160), .B2(n25070), .C1(n12162), .C2(n25569), .A(
        n12354), .ZN(n12351) );
  AOI221_X2 U4588 ( .B1(n12170), .B2(n25069), .C1(n12172), .C2(n25568), .A(
        n12359), .ZN(n12350) );
  OAI22_X2 U4589 ( .A1(n19192), .A2(n12175), .B1(n19166), .B2(n12176), .ZN(
        n12359) );
  AOI221_X2 U4592 ( .B1(n19173), .B2(n12177), .C1(n19164), .C2(n12178), .A(
        n12360), .ZN(n12349) );
  AOI221_X2 U4594 ( .B1(n19172), .B2(n12185), .C1(n19163), .C2(n12186), .A(
        n12363), .ZN(n12348) );
  OAI22_X2 U4595 ( .A1(n12188), .A2(n27953), .B1(n12190), .B2(n27873), .ZN(
        n12363) );
  NAND4_X2 U4596 ( .A1(n12366), .A2(n12367), .A3(n12368), .A4(n12369), .ZN(
        n12346) );
  AOI221_X2 U4597 ( .B1(n19195), .B2(n12196), .C1(n19194), .C2(n12197), .A(
        n12370), .ZN(n12369) );
  AOI221_X2 U4599 ( .B1(n12203), .B2(n25715), .C1(n12205), .C2(n25228), .A(
        n12374), .ZN(n12368) );
  OAI22_X2 U4600 ( .A1(n12208), .A2(n27905), .B1(n12210), .B2(n27921), .ZN(
        n12374) );
  AOI221_X2 U4603 ( .B1(n19178), .B2(n12212), .C1(n19177), .C2(n12213), .A(
        n12377), .ZN(n12367) );
  AOI221_X2 U4605 ( .B1(n12219), .B2(n25714), .C1(n12221), .C2(n25227), .A(
        n12381), .ZN(n12366) );
  OAI22_X2 U4606 ( .A1(n12224), .A2(n28065), .B1(n12226), .B2(n28081), .ZN(
        n12381) );
  NAND4_X2 U4611 ( .A1(n12387), .A2(n12388), .A3(n12389), .A4(n12390), .ZN(
        n12386) );
  AOI221_X2 U4612 ( .B1(n12160), .B2(n25068), .C1(n12162), .C2(n25567), .A(
        n12393), .ZN(n12390) );
  AOI221_X2 U4616 ( .B1(n12170), .B2(n25067), .C1(n12172), .C2(n25566), .A(
        n12398), .ZN(n12389) );
  OAI22_X2 U4617 ( .A1(n19155), .A2(n12175), .B1(n19129), .B2(n12176), .ZN(
        n12398) );
  AOI221_X2 U4620 ( .B1(n19136), .B2(n12177), .C1(n19127), .C2(n12178), .A(
        n12399), .ZN(n12388) );
  AOI221_X2 U4622 ( .B1(n19135), .B2(n12185), .C1(n19126), .C2(n12186), .A(
        n12402), .ZN(n12387) );
  OAI22_X2 U4623 ( .A1(n12188), .A2(n27952), .B1(n12190), .B2(n27872), .ZN(
        n12402) );
  NAND4_X2 U4624 ( .A1(n12405), .A2(n12406), .A3(n12407), .A4(n12408), .ZN(
        n12385) );
  AOI221_X2 U4625 ( .B1(n19158), .B2(n12196), .C1(n19157), .C2(n12197), .A(
        n12409), .ZN(n12408) );
  AOI221_X2 U4627 ( .B1(n12203), .B2(n25713), .C1(n12205), .C2(n25226), .A(
        n12413), .ZN(n12407) );
  OAI22_X2 U4628 ( .A1(n12208), .A2(n27904), .B1(n12210), .B2(n27920), .ZN(
        n12413) );
  AOI221_X2 U4631 ( .B1(n19141), .B2(n12212), .C1(n19140), .C2(n12213), .A(
        n12416), .ZN(n12406) );
  AOI221_X2 U4633 ( .B1(n12219), .B2(n25712), .C1(n12221), .C2(n25225), .A(
        n12420), .ZN(n12405) );
  OAI22_X2 U4634 ( .A1(n12224), .A2(n28064), .B1(n12226), .B2(n28080), .ZN(
        n12420) );
  NAND4_X2 U4639 ( .A1(n12426), .A2(n12427), .A3(n12428), .A4(n12429), .ZN(
        n12425) );
  AOI221_X2 U4640 ( .B1(n12160), .B2(n25066), .C1(n12162), .C2(n25565), .A(
        n12432), .ZN(n12429) );
  AOI221_X2 U4644 ( .B1(n12170), .B2(n25065), .C1(n12172), .C2(n25564), .A(
        n12437), .ZN(n12428) );
  OAI22_X2 U4645 ( .A1(n19118), .A2(n12175), .B1(n19092), .B2(n12176), .ZN(
        n12437) );
  AOI221_X2 U4648 ( .B1(n19099), .B2(n12177), .C1(n19090), .C2(n12178), .A(
        n12438), .ZN(n12427) );
  AOI221_X2 U4650 ( .B1(n19098), .B2(n12185), .C1(n19089), .C2(n12186), .A(
        n12441), .ZN(n12426) );
  OAI22_X2 U4651 ( .A1(n12188), .A2(n27951), .B1(n12190), .B2(n27871), .ZN(
        n12441) );
  NAND4_X2 U4652 ( .A1(n12444), .A2(n12445), .A3(n12446), .A4(n12447), .ZN(
        n12424) );
  AOI221_X2 U4653 ( .B1(n19121), .B2(n12196), .C1(n19120), .C2(n12197), .A(
        n12448), .ZN(n12447) );
  AOI221_X2 U4655 ( .B1(n12203), .B2(n25711), .C1(n12205), .C2(n25224), .A(
        n12452), .ZN(n12446) );
  OAI22_X2 U4656 ( .A1(n12208), .A2(n27903), .B1(n12210), .B2(n27919), .ZN(
        n12452) );
  AOI221_X2 U4659 ( .B1(n19104), .B2(n12212), .C1(n19103), .C2(n12213), .A(
        n12455), .ZN(n12445) );
  AOI221_X2 U4661 ( .B1(n12219), .B2(n25710), .C1(n12221), .C2(n25223), .A(
        n12459), .ZN(n12444) );
  OAI22_X2 U4662 ( .A1(n12224), .A2(n28063), .B1(n12226), .B2(n28079), .ZN(
        n12459) );
  NAND4_X2 U4667 ( .A1(n12465), .A2(n12466), .A3(n12467), .A4(n12468), .ZN(
        n12464) );
  AOI221_X2 U4668 ( .B1(n12160), .B2(n25064), .C1(n12162), .C2(n25563), .A(
        n12471), .ZN(n12468) );
  AOI221_X2 U4672 ( .B1(n12170), .B2(n25063), .C1(n12172), .C2(n25562), .A(
        n12476), .ZN(n12467) );
  OAI22_X2 U4673 ( .A1(n19081), .A2(n12175), .B1(n19055), .B2(n12176), .ZN(
        n12476) );
  AOI221_X2 U4676 ( .B1(n19062), .B2(n12177), .C1(n19053), .C2(n12178), .A(
        n12477), .ZN(n12466) );
  AOI221_X2 U4678 ( .B1(n19061), .B2(n12185), .C1(n19052), .C2(n12186), .A(
        n12480), .ZN(n12465) );
  OAI22_X2 U4679 ( .A1(n12188), .A2(n27950), .B1(n12190), .B2(n27870), .ZN(
        n12480) );
  NAND4_X2 U4680 ( .A1(n12483), .A2(n12484), .A3(n12485), .A4(n12486), .ZN(
        n12463) );
  AOI221_X2 U4681 ( .B1(n19084), .B2(n12196), .C1(n19083), .C2(n12197), .A(
        n12487), .ZN(n12486) );
  AOI221_X2 U4683 ( .B1(n12203), .B2(n25709), .C1(n12205), .C2(n25222), .A(
        n12491), .ZN(n12485) );
  OAI22_X2 U4684 ( .A1(n12208), .A2(n27902), .B1(n12210), .B2(n27918), .ZN(
        n12491) );
  AOI221_X2 U4687 ( .B1(n19067), .B2(n12212), .C1(n19066), .C2(n12213), .A(
        n12494), .ZN(n12484) );
  AOI221_X2 U4689 ( .B1(n12219), .B2(n25708), .C1(n12221), .C2(n25221), .A(
        n12498), .ZN(n12483) );
  OAI22_X2 U4690 ( .A1(n12224), .A2(n28062), .B1(n12226), .B2(n28078), .ZN(
        n12498) );
  NAND4_X2 U4695 ( .A1(n12504), .A2(n12505), .A3(n12506), .A4(n12507), .ZN(
        n12503) );
  AOI221_X2 U4696 ( .B1(n12160), .B2(n25277), .C1(n12162), .C2(n24910), .A(
        n12510), .ZN(n12507) );
  AOI221_X2 U4700 ( .B1(n12170), .B2(n25276), .C1(n12172), .C2(n24909), .A(
        n12515), .ZN(n12506) );
  OAI22_X2 U4701 ( .A1(n19044), .A2(n12175), .B1(n19018), .B2(n12176), .ZN(
        n12515) );
  AOI221_X2 U4704 ( .B1(n19025), .B2(n12177), .C1(n19016), .C2(n12178), .A(
        n12516), .ZN(n12505) );
  AOI221_X2 U4706 ( .B1(n19024), .B2(n12185), .C1(n19015), .C2(n12186), .A(
        n12519), .ZN(n12504) );
  OAI22_X2 U4707 ( .A1(n12188), .A2(n27949), .B1(n12190), .B2(n27869), .ZN(
        n12519) );
  NAND4_X2 U4708 ( .A1(n12522), .A2(n12523), .A3(n12524), .A4(n12525), .ZN(
        n12502) );
  AOI221_X2 U4709 ( .B1(n19047), .B2(n12196), .C1(n19046), .C2(n12197), .A(
        n12526), .ZN(n12525) );
  AOI221_X2 U4711 ( .B1(n12203), .B2(n25275), .C1(n12205), .C2(n24908), .A(
        n12530), .ZN(n12524) );
  OAI22_X2 U4712 ( .A1(n12208), .A2(n27901), .B1(n12210), .B2(n27917), .ZN(
        n12530) );
  AOI221_X2 U4715 ( .B1(n19030), .B2(n12212), .C1(n19029), .C2(n12213), .A(
        n12533), .ZN(n12523) );
  AOI221_X2 U4717 ( .B1(n12219), .B2(n25274), .C1(n12221), .C2(n24907), .A(
        n12537), .ZN(n12522) );
  OAI22_X2 U4718 ( .A1(n12224), .A2(n28061), .B1(n12226), .B2(n28077), .ZN(
        n12537) );
  NAND4_X2 U4723 ( .A1(n12543), .A2(n12544), .A3(n12545), .A4(n12546), .ZN(
        n12542) );
  AOI221_X2 U4724 ( .B1(n12160), .B2(n25062), .C1(n12162), .C2(n25561), .A(
        n12549), .ZN(n12546) );
  AOI221_X2 U4728 ( .B1(n12170), .B2(n25061), .C1(n12172), .C2(n25560), .A(
        n12554), .ZN(n12545) );
  OAI22_X2 U4729 ( .A1(n19007), .A2(n12175), .B1(n18981), .B2(n12176), .ZN(
        n12554) );
  AOI221_X2 U4732 ( .B1(n18988), .B2(n12177), .C1(n18979), .C2(n12178), .A(
        n12555), .ZN(n12544) );
  AOI221_X2 U4734 ( .B1(n18987), .B2(n12185), .C1(n18978), .C2(n12186), .A(
        n12558), .ZN(n12543) );
  OAI22_X2 U4735 ( .A1(n12188), .A2(n27948), .B1(n12190), .B2(n27868), .ZN(
        n12558) );
  NAND4_X2 U4736 ( .A1(n12561), .A2(n12562), .A3(n12563), .A4(n12564), .ZN(
        n12541) );
  AOI221_X2 U4737 ( .B1(n19010), .B2(n12196), .C1(n19009), .C2(n12197), .A(
        n12565), .ZN(n12564) );
  AOI221_X2 U4739 ( .B1(n12203), .B2(n25707), .C1(n12205), .C2(n25220), .A(
        n12569), .ZN(n12563) );
  OAI22_X2 U4740 ( .A1(n12208), .A2(n27900), .B1(n12210), .B2(n27916), .ZN(
        n12569) );
  AOI221_X2 U4743 ( .B1(n18993), .B2(n12212), .C1(n18992), .C2(n12213), .A(
        n12572), .ZN(n12562) );
  AOI221_X2 U4745 ( .B1(n12219), .B2(n25706), .C1(n12221), .C2(n25219), .A(
        n12576), .ZN(n12561) );
  OAI22_X2 U4746 ( .A1(n12224), .A2(n28060), .B1(n12226), .B2(n28076), .ZN(
        n12576) );
  NAND4_X2 U4751 ( .A1(n12582), .A2(n12583), .A3(n12584), .A4(n12585), .ZN(
        n12581) );
  AOI221_X2 U4752 ( .B1(n12160), .B2(n25060), .C1(n12162), .C2(n25559), .A(
        n12588), .ZN(n12585) );
  AOI221_X2 U4756 ( .B1(n12170), .B2(n25059), .C1(n12172), .C2(n25558), .A(
        n12593), .ZN(n12584) );
  OAI22_X2 U4757 ( .A1(n18970), .A2(n12175), .B1(n18944), .B2(n12176), .ZN(
        n12593) );
  AOI221_X2 U4760 ( .B1(n18951), .B2(n12177), .C1(n18942), .C2(n12178), .A(
        n12594), .ZN(n12583) );
  AOI221_X2 U4762 ( .B1(n18950), .B2(n12185), .C1(n18941), .C2(n12186), .A(
        n12597), .ZN(n12582) );
  OAI22_X2 U4763 ( .A1(n12188), .A2(n27947), .B1(n12190), .B2(n27867), .ZN(
        n12597) );
  NAND4_X2 U4764 ( .A1(n12600), .A2(n12601), .A3(n12602), .A4(n12603), .ZN(
        n12580) );
  AOI221_X2 U4765 ( .B1(n18973), .B2(n12196), .C1(n18972), .C2(n12197), .A(
        n12604), .ZN(n12603) );
  AOI221_X2 U4767 ( .B1(n12203), .B2(n25705), .C1(n12205), .C2(n25218), .A(
        n12608), .ZN(n12602) );
  OAI22_X2 U4768 ( .A1(n12208), .A2(n27899), .B1(n12210), .B2(n27915), .ZN(
        n12608) );
  AOI221_X2 U4771 ( .B1(n18956), .B2(n12212), .C1(n18955), .C2(n12213), .A(
        n12611), .ZN(n12601) );
  AOI221_X2 U4773 ( .B1(n12219), .B2(n25704), .C1(n12221), .C2(n25217), .A(
        n12615), .ZN(n12600) );
  OAI22_X2 U4774 ( .A1(n12224), .A2(n28059), .B1(n12226), .B2(n28075), .ZN(
        n12615) );
  NAND4_X2 U4779 ( .A1(n12621), .A2(n12622), .A3(n12623), .A4(n12624), .ZN(
        n12620) );
  AOI221_X2 U4780 ( .B1(n12160), .B2(n25058), .C1(n12162), .C2(n25557), .A(
        n12627), .ZN(n12624) );
  AOI221_X2 U4784 ( .B1(n12170), .B2(n25057), .C1(n12172), .C2(n25556), .A(
        n12632), .ZN(n12623) );
  OAI22_X2 U4785 ( .A1(n18933), .A2(n12175), .B1(n18907), .B2(n12176), .ZN(
        n12632) );
  AOI221_X2 U4788 ( .B1(n18914), .B2(n12177), .C1(n18905), .C2(n12178), .A(
        n12633), .ZN(n12622) );
  AOI221_X2 U4790 ( .B1(n18913), .B2(n12185), .C1(n18904), .C2(n12186), .A(
        n12636), .ZN(n12621) );
  OAI22_X2 U4791 ( .A1(n12188), .A2(n27946), .B1(n12190), .B2(n27866), .ZN(
        n12636) );
  NAND4_X2 U4792 ( .A1(n12639), .A2(n12640), .A3(n12641), .A4(n12642), .ZN(
        n12619) );
  AOI221_X2 U4793 ( .B1(n18936), .B2(n12196), .C1(n18935), .C2(n12197), .A(
        n12643), .ZN(n12642) );
  AOI221_X2 U4795 ( .B1(n12203), .B2(n25703), .C1(n12205), .C2(n25216), .A(
        n12647), .ZN(n12641) );
  OAI22_X2 U4796 ( .A1(n12208), .A2(n27898), .B1(n12210), .B2(n27914), .ZN(
        n12647) );
  AOI221_X2 U4799 ( .B1(n18919), .B2(n12212), .C1(n18918), .C2(n12213), .A(
        n12650), .ZN(n12640) );
  AOI221_X2 U4801 ( .B1(n12219), .B2(n25702), .C1(n12221), .C2(n25215), .A(
        n12654), .ZN(n12639) );
  OAI22_X2 U4802 ( .A1(n12224), .A2(n28058), .B1(n12226), .B2(n28074), .ZN(
        n12654) );
  NAND4_X2 U4807 ( .A1(n12660), .A2(n12661), .A3(n12662), .A4(n12663), .ZN(
        n12659) );
  AOI221_X2 U4808 ( .B1(n12160), .B2(n25273), .C1(n12162), .C2(n24906), .A(
        n12666), .ZN(n12663) );
  AOI221_X2 U4812 ( .B1(n12170), .B2(n25272), .C1(n12172), .C2(n24905), .A(
        n12671), .ZN(n12662) );
  OAI22_X2 U4813 ( .A1(n18896), .A2(n12175), .B1(n18870), .B2(n12176), .ZN(
        n12671) );
  AOI221_X2 U4816 ( .B1(n18877), .B2(n12177), .C1(n18868), .C2(n12178), .A(
        n12672), .ZN(n12661) );
  AOI221_X2 U4818 ( .B1(n18876), .B2(n12185), .C1(n18867), .C2(n12186), .A(
        n12675), .ZN(n12660) );
  OAI22_X2 U4819 ( .A1(n12188), .A2(n27945), .B1(n12190), .B2(n27865), .ZN(
        n12675) );
  NAND4_X2 U4820 ( .A1(n12678), .A2(n12679), .A3(n12680), .A4(n12681), .ZN(
        n12658) );
  AOI221_X2 U4821 ( .B1(n18899), .B2(n12196), .C1(n18898), .C2(n12197), .A(
        n12682), .ZN(n12681) );
  AOI221_X2 U4823 ( .B1(n12203), .B2(n25271), .C1(n12205), .C2(n24904), .A(
        n12686), .ZN(n12680) );
  OAI22_X2 U4824 ( .A1(n12208), .A2(n27897), .B1(n12210), .B2(n27913), .ZN(
        n12686) );
  AOI221_X2 U4827 ( .B1(n18882), .B2(n12212), .C1(n18881), .C2(n12213), .A(
        n12689), .ZN(n12679) );
  AOI221_X2 U4829 ( .B1(n12219), .B2(n25270), .C1(n12221), .C2(n24903), .A(
        n12693), .ZN(n12678) );
  OAI22_X2 U4830 ( .A1(n12224), .A2(n28057), .B1(n12226), .B2(n28073), .ZN(
        n12693) );
  NAND4_X2 U4835 ( .A1(n12699), .A2(n12700), .A3(n12701), .A4(n12702), .ZN(
        n12698) );
  AOI221_X2 U4836 ( .B1(n12160), .B2(n25056), .C1(n12162), .C2(n25555), .A(
        n12705), .ZN(n12702) );
  AOI221_X2 U4840 ( .B1(n12170), .B2(n25055), .C1(n12172), .C2(n25554), .A(
        n12710), .ZN(n12701) );
  OAI22_X2 U4841 ( .A1(n18859), .A2(n12175), .B1(n18833), .B2(n12176), .ZN(
        n12710) );
  AOI221_X2 U4844 ( .B1(n18840), .B2(n12177), .C1(n18831), .C2(n12178), .A(
        n12711), .ZN(n12700) );
  AOI221_X2 U4846 ( .B1(n18839), .B2(n12185), .C1(n18830), .C2(n12186), .A(
        n12714), .ZN(n12699) );
  OAI22_X2 U4847 ( .A1(n12188), .A2(n27944), .B1(n12190), .B2(n27864), .ZN(
        n12714) );
  NAND4_X2 U4848 ( .A1(n12717), .A2(n12718), .A3(n12719), .A4(n12720), .ZN(
        n12697) );
  AOI221_X2 U4849 ( .B1(n18862), .B2(n12196), .C1(n18861), .C2(n12197), .A(
        n12721), .ZN(n12720) );
  AOI221_X2 U4851 ( .B1(n12203), .B2(n25701), .C1(n12205), .C2(n25214), .A(
        n12725), .ZN(n12719) );
  OAI22_X2 U4852 ( .A1(n12208), .A2(n27896), .B1(n12210), .B2(n27912), .ZN(
        n12725) );
  AOI221_X2 U4855 ( .B1(n18845), .B2(n12212), .C1(n18844), .C2(n12213), .A(
        n12728), .ZN(n12718) );
  AOI221_X2 U4857 ( .B1(n12219), .B2(n25700), .C1(n12221), .C2(n25213), .A(
        n12732), .ZN(n12717) );
  OAI22_X2 U4858 ( .A1(n12224), .A2(n28056), .B1(n12226), .B2(n28072), .ZN(
        n12732) );
  NAND4_X2 U4863 ( .A1(n12738), .A2(n12739), .A3(n12740), .A4(n12741), .ZN(
        n12737) );
  AOI221_X2 U4864 ( .B1(n12160), .B2(n25269), .C1(n12162), .C2(n24902), .A(
        n12744), .ZN(n12741) );
  AOI221_X2 U4868 ( .B1(n12170), .B2(n25268), .C1(n12172), .C2(n24901), .A(
        n12749), .ZN(n12740) );
  OAI22_X2 U4869 ( .A1(n18822), .A2(n12175), .B1(n18796), .B2(n12176), .ZN(
        n12749) );
  AOI221_X2 U4872 ( .B1(n18803), .B2(n12177), .C1(n18794), .C2(n12178), .A(
        n12750), .ZN(n12739) );
  AOI221_X2 U4874 ( .B1(n18802), .B2(n12185), .C1(n18793), .C2(n12186), .A(
        n12753), .ZN(n12738) );
  OAI22_X2 U4875 ( .A1(n12188), .A2(n27943), .B1(n12190), .B2(n27863), .ZN(
        n12753) );
  NAND4_X2 U4876 ( .A1(n12756), .A2(n12757), .A3(n12758), .A4(n12759), .ZN(
        n12736) );
  AOI221_X2 U4877 ( .B1(n18825), .B2(n12196), .C1(n18824), .C2(n12197), .A(
        n12760), .ZN(n12759) );
  AOI221_X2 U4879 ( .B1(n12203), .B2(n25267), .C1(n12205), .C2(n24900), .A(
        n12764), .ZN(n12758) );
  OAI22_X2 U4880 ( .A1(n12208), .A2(n27895), .B1(n12210), .B2(n27911), .ZN(
        n12764) );
  AOI221_X2 U4883 ( .B1(n18808), .B2(n12212), .C1(n18807), .C2(n12213), .A(
        n12767), .ZN(n12757) );
  AOI221_X2 U4885 ( .B1(n12219), .B2(n25266), .C1(n12221), .C2(n24899), .A(
        n12771), .ZN(n12756) );
  OAI22_X2 U4886 ( .A1(n12224), .A2(n28055), .B1(n12226), .B2(n28071), .ZN(
        n12771) );
  NAND4_X2 U4891 ( .A1(n12777), .A2(n12778), .A3(n12779), .A4(n12780), .ZN(
        n12776) );
  AOI221_X2 U4892 ( .B1(n12160), .B2(n25054), .C1(n12162), .C2(n25553), .A(
        n12783), .ZN(n12780) );
  AOI221_X2 U4901 ( .B1(n12170), .B2(n25053), .C1(n12172), .C2(n25552), .A(
        n12794), .ZN(n12779) );
  OAI22_X2 U4902 ( .A1(n18785), .A2(n12175), .B1(n18759), .B2(n12176), .ZN(
        n12794) );
  AOI221_X2 U4909 ( .B1(n18766), .B2(n12177), .C1(n18757), .C2(n12178), .A(
        n12796), .ZN(n12778) );
  AOI221_X2 U4916 ( .B1(n18765), .B2(n12185), .C1(n18756), .C2(n12186), .A(
        n12800), .ZN(n12777) );
  OAI22_X2 U4917 ( .A1(n12188), .A2(n27942), .B1(n12190), .B2(n27862), .ZN(
        n12800) );
  NAND4_X2 U4922 ( .A1(n12804), .A2(n12805), .A3(n12806), .A4(n12807), .ZN(
        n12775) );
  AOI221_X2 U4923 ( .B1(n18788), .B2(n12196), .C1(n18787), .C2(n12197), .A(
        n12808), .ZN(n12807) );
  AOI221_X2 U4931 ( .B1(n12203), .B2(n25699), .C1(n12205), .C2(n25212), .A(
        n12820), .ZN(n12806) );
  OAI22_X2 U4932 ( .A1(n12208), .A2(n27894), .B1(n12210), .B2(n27910), .ZN(
        n12820) );
  AOI221_X2 U4939 ( .B1(n18771), .B2(n12212), .C1(n18770), .C2(n12213), .A(
        n12823), .ZN(n12805) );
  AOI221_X2 U4948 ( .B1(n12219), .B2(n25698), .C1(n12221), .C2(n25211), .A(
        n12835), .ZN(n12804) );
  OAI22_X2 U4949 ( .A1(n12224), .A2(n28054), .B1(n12226), .B2(n28070), .ZN(
        n12835) );
  OAI22_X2 U4957 ( .A1(n26337), .A2(n28054), .B1(n26134), .B2(n12843), .ZN(
        n23104) );
  OAI22_X2 U4959 ( .A1(n26337), .A2(n28055), .B1(n26133), .B2(n12843), .ZN(
        n23105) );
  OAI22_X2 U4961 ( .A1(n26337), .A2(n28056), .B1(n26132), .B2(n12843), .ZN(
        n23106) );
  OAI22_X2 U4963 ( .A1(n26337), .A2(n28057), .B1(n26131), .B2(n12843), .ZN(
        n23107) );
  OAI22_X2 U4965 ( .A1(n26337), .A2(n28058), .B1(n26279), .B2(n12843), .ZN(
        n23108) );
  OAI22_X2 U4967 ( .A1(n26337), .A2(n28059), .B1(n26278), .B2(n12843), .ZN(
        n23109) );
  OAI22_X2 U4969 ( .A1(n26337), .A2(n28060), .B1(n26277), .B2(n12843), .ZN(
        n23110) );
  OAI22_X2 U4971 ( .A1(n26337), .A2(n28061), .B1(n26276), .B2(n12843), .ZN(
        n23111) );
  OAI22_X2 U4973 ( .A1(n26337), .A2(n28062), .B1(n26275), .B2(n12843), .ZN(
        n23112) );
  OAI22_X2 U4975 ( .A1(n26337), .A2(n28063), .B1(n26274), .B2(n12843), .ZN(
        n23113) );
  OAI22_X2 U4977 ( .A1(n26337), .A2(n28064), .B1(n26273), .B2(n12843), .ZN(
        n23114) );
  OAI22_X2 U4979 ( .A1(n26337), .A2(n28065), .B1(n26272), .B2(n12843), .ZN(
        n23115) );
  OAI22_X2 U4981 ( .A1(n26337), .A2(n28066), .B1(n26271), .B2(n12843), .ZN(
        n23116) );
  OAI22_X2 U4983 ( .A1(n26337), .A2(n28067), .B1(n26270), .B2(n12843), .ZN(
        n23117) );
  OAI22_X2 U4985 ( .A1(n26337), .A2(n28068), .B1(n26269), .B2(n12843), .ZN(
        n23118) );
  OAI22_X2 U4987 ( .A1(n26337), .A2(n28069), .B1(n26268), .B2(n12843), .ZN(
        n23119) );
  OAI22_X2 U4991 ( .A1(n26336), .A2(n28070), .B1(n26134), .B2(n12846), .ZN(
        n23120) );
  OAI22_X2 U4993 ( .A1(n26336), .A2(n28071), .B1(n26133), .B2(n12846), .ZN(
        n23121) );
  OAI22_X2 U4995 ( .A1(n26336), .A2(n28072), .B1(n26132), .B2(n12846), .ZN(
        n23122) );
  OAI22_X2 U4997 ( .A1(n26336), .A2(n28073), .B1(n26131), .B2(n12846), .ZN(
        n23123) );
  OAI22_X2 U4999 ( .A1(n26336), .A2(n28074), .B1(n26279), .B2(n12846), .ZN(
        n23124) );
  OAI22_X2 U5001 ( .A1(n26336), .A2(n28075), .B1(n26278), .B2(n12846), .ZN(
        n23125) );
  OAI22_X2 U5003 ( .A1(n26336), .A2(n28076), .B1(n26277), .B2(n12846), .ZN(
        n23126) );
  OAI22_X2 U5005 ( .A1(n26336), .A2(n28077), .B1(n26276), .B2(n12846), .ZN(
        n23127) );
  OAI22_X2 U5007 ( .A1(n26336), .A2(n28078), .B1(n26275), .B2(n12846), .ZN(
        n23128) );
  OAI22_X2 U5009 ( .A1(n26336), .A2(n28079), .B1(n26274), .B2(n12846), .ZN(
        n23129) );
  OAI22_X2 U5011 ( .A1(n26336), .A2(n28080), .B1(n26273), .B2(n12846), .ZN(
        n23130) );
  OAI22_X2 U5013 ( .A1(n26336), .A2(n28081), .B1(n26272), .B2(n12846), .ZN(
        n23131) );
  OAI22_X2 U5015 ( .A1(n26336), .A2(n28082), .B1(n26271), .B2(n12846), .ZN(
        n23132) );
  OAI22_X2 U5017 ( .A1(n26336), .A2(n28083), .B1(n26270), .B2(n12846), .ZN(
        n23133) );
  OAI22_X2 U5019 ( .A1(n26336), .A2(n28084), .B1(n26269), .B2(n12846), .ZN(
        n23134) );
  OAI22_X2 U5021 ( .A1(n26336), .A2(n28085), .B1(n26268), .B2(n12846), .ZN(
        n23135) );
  OAI22_X2 U5025 ( .A1(n26335), .A2(n28086), .B1(n26134), .B2(n12849), .ZN(
        n23136) );
  OAI22_X2 U5027 ( .A1(n26335), .A2(n28087), .B1(n26133), .B2(n12849), .ZN(
        n23137) );
  OAI22_X2 U5029 ( .A1(n26335), .A2(n28088), .B1(n26132), .B2(n12849), .ZN(
        n23138) );
  OAI22_X2 U5031 ( .A1(n26335), .A2(n28089), .B1(n26131), .B2(n12849), .ZN(
        n23139) );
  OAI22_X2 U5033 ( .A1(n26335), .A2(n28090), .B1(n26279), .B2(n12849), .ZN(
        n23140) );
  OAI22_X2 U5035 ( .A1(n26335), .A2(n28091), .B1(n26278), .B2(n12849), .ZN(
        n23141) );
  OAI22_X2 U5037 ( .A1(n26335), .A2(n28092), .B1(n26277), .B2(n12849), .ZN(
        n23142) );
  OAI22_X2 U5039 ( .A1(n26335), .A2(n28093), .B1(n26276), .B2(n12849), .ZN(
        n23143) );
  OAI22_X2 U5041 ( .A1(n26335), .A2(n28094), .B1(n26275), .B2(n12849), .ZN(
        n23144) );
  OAI22_X2 U5043 ( .A1(n26335), .A2(n28095), .B1(n26274), .B2(n12849), .ZN(
        n23145) );
  OAI22_X2 U5045 ( .A1(n26335), .A2(n28096), .B1(n26273), .B2(n12849), .ZN(
        n23146) );
  OAI22_X2 U5047 ( .A1(n26335), .A2(n28097), .B1(n26272), .B2(n12849), .ZN(
        n23147) );
  OAI22_X2 U5049 ( .A1(n26335), .A2(n28098), .B1(n26271), .B2(n12849), .ZN(
        n23148) );
  OAI22_X2 U5051 ( .A1(n26335), .A2(n28099), .B1(n26270), .B2(n12849), .ZN(
        n23149) );
  OAI22_X2 U5053 ( .A1(n26335), .A2(n28100), .B1(n26269), .B2(n12849), .ZN(
        n23150) );
  OAI22_X2 U5055 ( .A1(n26335), .A2(n28101), .B1(n26268), .B2(n12849), .ZN(
        n23151) );
  OAI22_X2 U5059 ( .A1(n26334), .A2(n28102), .B1(n26134), .B2(n12853), .ZN(
        n23152) );
  OAI22_X2 U5061 ( .A1(n26334), .A2(n28103), .B1(n26133), .B2(n12853), .ZN(
        n23153) );
  OAI22_X2 U5063 ( .A1(n26334), .A2(n28104), .B1(n26132), .B2(n12853), .ZN(
        n23154) );
  OAI22_X2 U5065 ( .A1(n26334), .A2(n28105), .B1(n26131), .B2(n12853), .ZN(
        n23155) );
  OAI22_X2 U5067 ( .A1(n26334), .A2(n28106), .B1(n26279), .B2(n12853), .ZN(
        n23156) );
  OAI22_X2 U5069 ( .A1(n26334), .A2(n28107), .B1(n26278), .B2(n12853), .ZN(
        n23157) );
  OAI22_X2 U5071 ( .A1(n26334), .A2(n28108), .B1(n26277), .B2(n12853), .ZN(
        n23158) );
  OAI22_X2 U5073 ( .A1(n26334), .A2(n28109), .B1(n26276), .B2(n12853), .ZN(
        n23159) );
  OAI22_X2 U5075 ( .A1(n26334), .A2(n28110), .B1(n26275), .B2(n12853), .ZN(
        n23160) );
  OAI22_X2 U5077 ( .A1(n26334), .A2(n28111), .B1(n26274), .B2(n12853), .ZN(
        n23161) );
  OAI22_X2 U5079 ( .A1(n26334), .A2(n28112), .B1(n26273), .B2(n12853), .ZN(
        n23162) );
  OAI22_X2 U5081 ( .A1(n26334), .A2(n28113), .B1(n26272), .B2(n12853), .ZN(
        n23163) );
  OAI22_X2 U5083 ( .A1(n26334), .A2(n28114), .B1(n26271), .B2(n12853), .ZN(
        n23164) );
  OAI22_X2 U5085 ( .A1(n26334), .A2(n28115), .B1(n26270), .B2(n12853), .ZN(
        n23165) );
  OAI22_X2 U5087 ( .A1(n26334), .A2(n28116), .B1(n26269), .B2(n12853), .ZN(
        n23166) );
  OAI22_X2 U5089 ( .A1(n26334), .A2(n28117), .B1(n26268), .B2(n12853), .ZN(
        n23167) );
  OAI22_X2 U5093 ( .A1(n26333), .A2(n28118), .B1(n26134), .B2(n12872), .ZN(
        n23168) );
  OAI22_X2 U5095 ( .A1(n26333), .A2(n28119), .B1(n26133), .B2(n12872), .ZN(
        n23169) );
  OAI22_X2 U5097 ( .A1(n26333), .A2(n28120), .B1(n26132), .B2(n12872), .ZN(
        n23170) );
  OAI22_X2 U5099 ( .A1(n26333), .A2(n28121), .B1(n26131), .B2(n12872), .ZN(
        n23171) );
  OAI22_X2 U5101 ( .A1(n26333), .A2(n28122), .B1(n26279), .B2(n12872), .ZN(
        n23172) );
  OAI22_X2 U5103 ( .A1(n26333), .A2(n28123), .B1(n26278), .B2(n12872), .ZN(
        n23173) );
  OAI22_X2 U5105 ( .A1(n26333), .A2(n28124), .B1(n26277), .B2(n12872), .ZN(
        n23174) );
  OAI22_X2 U5107 ( .A1(n26333), .A2(n28125), .B1(n26276), .B2(n12872), .ZN(
        n23175) );
  OAI22_X2 U5109 ( .A1(n26333), .A2(n28126), .B1(n26275), .B2(n12872), .ZN(
        n23176) );
  OAI22_X2 U5111 ( .A1(n26333), .A2(n28127), .B1(n26274), .B2(n12872), .ZN(
        n23177) );
  OAI22_X2 U5113 ( .A1(n26333), .A2(n28128), .B1(n26273), .B2(n12872), .ZN(
        n23178) );
  OAI22_X2 U5115 ( .A1(n26333), .A2(n28129), .B1(n26272), .B2(n12872), .ZN(
        n23179) );
  OAI22_X2 U5117 ( .A1(n26333), .A2(n28130), .B1(n26271), .B2(n12872), .ZN(
        n23180) );
  OAI22_X2 U5119 ( .A1(n26333), .A2(n28131), .B1(n26270), .B2(n12872), .ZN(
        n23181) );
  OAI22_X2 U5121 ( .A1(n26333), .A2(n28132), .B1(n26269), .B2(n12872), .ZN(
        n23182) );
  OAI22_X2 U5123 ( .A1(n26333), .A2(n28133), .B1(n26268), .B2(n12872), .ZN(
        n23183) );
  OAI22_X2 U5128 ( .A1(n26328), .A2(n27974), .B1(n26134), .B2(n12892), .ZN(
        n23184) );
  OAI22_X2 U5130 ( .A1(n26328), .A2(n27975), .B1(n26133), .B2(n12892), .ZN(
        n23185) );
  OAI22_X2 U5132 ( .A1(n26328), .A2(n27976), .B1(n26132), .B2(n12892), .ZN(
        n23186) );
  OAI22_X2 U5134 ( .A1(n26328), .A2(n27977), .B1(n26131), .B2(n12892), .ZN(
        n23187) );
  OAI22_X2 U5136 ( .A1(n26328), .A2(n27978), .B1(n26279), .B2(n12892), .ZN(
        n23188) );
  OAI22_X2 U5138 ( .A1(n26328), .A2(n27979), .B1(n26278), .B2(n12892), .ZN(
        n23189) );
  OAI22_X2 U5140 ( .A1(n26328), .A2(n27980), .B1(n26277), .B2(n12892), .ZN(
        n23190) );
  OAI22_X2 U5142 ( .A1(n26328), .A2(n27981), .B1(n26276), .B2(n12892), .ZN(
        n23191) );
  OAI22_X2 U5144 ( .A1(n26328), .A2(n27982), .B1(n26275), .B2(n12892), .ZN(
        n23192) );
  OAI22_X2 U5146 ( .A1(n26328), .A2(n27983), .B1(n26274), .B2(n12892), .ZN(
        n23193) );
  OAI22_X2 U5148 ( .A1(n26328), .A2(n27984), .B1(n26273), .B2(n12892), .ZN(
        n23194) );
  OAI22_X2 U5150 ( .A1(n26328), .A2(n27985), .B1(n26272), .B2(n12892), .ZN(
        n23195) );
  OAI22_X2 U5152 ( .A1(n26328), .A2(n27986), .B1(n26271), .B2(n12892), .ZN(
        n23196) );
  OAI22_X2 U5154 ( .A1(n26328), .A2(n27987), .B1(n26270), .B2(n12892), .ZN(
        n23197) );
  OAI22_X2 U5156 ( .A1(n26328), .A2(n27988), .B1(n26269), .B2(n12892), .ZN(
        n23198) );
  OAI22_X2 U5158 ( .A1(n26328), .A2(n27989), .B1(n26268), .B2(n12892), .ZN(
        n23199) );
  OAI22_X2 U5162 ( .A1(n26327), .A2(n27990), .B1(n26134), .B2(n12910), .ZN(
        n23200) );
  OAI22_X2 U5164 ( .A1(n26327), .A2(n27991), .B1(n26133), .B2(n12910), .ZN(
        n23201) );
  OAI22_X2 U5166 ( .A1(n26327), .A2(n27992), .B1(n26132), .B2(n12910), .ZN(
        n23202) );
  OAI22_X2 U5168 ( .A1(n26327), .A2(n27993), .B1(n26131), .B2(n12910), .ZN(
        n23203) );
  OAI22_X2 U5170 ( .A1(n26327), .A2(n27994), .B1(n26279), .B2(n12910), .ZN(
        n23204) );
  OAI22_X2 U5172 ( .A1(n26327), .A2(n27995), .B1(n26278), .B2(n12910), .ZN(
        n23205) );
  OAI22_X2 U5174 ( .A1(n26327), .A2(n27996), .B1(n26277), .B2(n12910), .ZN(
        n23206) );
  OAI22_X2 U5176 ( .A1(n26327), .A2(n27997), .B1(n26276), .B2(n12910), .ZN(
        n23207) );
  OAI22_X2 U5178 ( .A1(n26327), .A2(n27998), .B1(n26275), .B2(n12910), .ZN(
        n23208) );
  OAI22_X2 U5180 ( .A1(n26327), .A2(n27999), .B1(n26274), .B2(n12910), .ZN(
        n23209) );
  OAI22_X2 U5182 ( .A1(n26327), .A2(n28000), .B1(n26273), .B2(n12910), .ZN(
        n23210) );
  OAI22_X2 U5184 ( .A1(n26327), .A2(n28001), .B1(n26272), .B2(n12910), .ZN(
        n23211) );
  OAI22_X2 U5186 ( .A1(n26327), .A2(n28002), .B1(n26271), .B2(n12910), .ZN(
        n23212) );
  OAI22_X2 U5188 ( .A1(n26327), .A2(n28003), .B1(n26270), .B2(n12910), .ZN(
        n23213) );
  OAI22_X2 U5190 ( .A1(n26327), .A2(n28004), .B1(n26269), .B2(n12910), .ZN(
        n23214) );
  OAI22_X2 U5192 ( .A1(n26327), .A2(n28005), .B1(n26268), .B2(n12910), .ZN(
        n23215) );
  OAI22_X2 U5196 ( .A1(n26326), .A2(n28006), .B1(n26134), .B2(n12927), .ZN(
        n23216) );
  OAI22_X2 U5198 ( .A1(n26326), .A2(n28007), .B1(n26133), .B2(n12927), .ZN(
        n23217) );
  OAI22_X2 U5200 ( .A1(n26326), .A2(n28008), .B1(n26132), .B2(n12927), .ZN(
        n23218) );
  OAI22_X2 U5202 ( .A1(n26326), .A2(n28009), .B1(n26131), .B2(n12927), .ZN(
        n23219) );
  OAI22_X2 U5204 ( .A1(n26326), .A2(n28010), .B1(n26279), .B2(n12927), .ZN(
        n23220) );
  OAI22_X2 U5206 ( .A1(n26326), .A2(n28011), .B1(n26278), .B2(n12927), .ZN(
        n23221) );
  OAI22_X2 U5208 ( .A1(n26326), .A2(n28012), .B1(n26277), .B2(n12927), .ZN(
        n23222) );
  OAI22_X2 U5210 ( .A1(n26326), .A2(n28013), .B1(n26276), .B2(n12927), .ZN(
        n23223) );
  OAI22_X2 U5212 ( .A1(n26326), .A2(n28014), .B1(n26275), .B2(n12927), .ZN(
        n23224) );
  OAI22_X2 U5214 ( .A1(n26326), .A2(n28015), .B1(n26274), .B2(n12927), .ZN(
        n23225) );
  OAI22_X2 U5216 ( .A1(n26326), .A2(n28016), .B1(n26273), .B2(n12927), .ZN(
        n23226) );
  OAI22_X2 U5218 ( .A1(n26326), .A2(n28017), .B1(n26272), .B2(n12927), .ZN(
        n23227) );
  OAI22_X2 U5220 ( .A1(n26326), .A2(n28018), .B1(n26271), .B2(n12927), .ZN(
        n23228) );
  OAI22_X2 U5222 ( .A1(n26326), .A2(n28019), .B1(n26270), .B2(n12927), .ZN(
        n23229) );
  OAI22_X2 U5224 ( .A1(n26326), .A2(n28020), .B1(n26269), .B2(n12927), .ZN(
        n23230) );
  OAI22_X2 U5226 ( .A1(n26326), .A2(n28021), .B1(n26268), .B2(n12927), .ZN(
        n23231) );
  OAI22_X2 U5230 ( .A1(n26325), .A2(n28022), .B1(n26134), .B2(n12930), .ZN(
        n23232) );
  OAI22_X2 U5232 ( .A1(n26325), .A2(n28023), .B1(n26133), .B2(n12930), .ZN(
        n23233) );
  OAI22_X2 U5234 ( .A1(n26325), .A2(n28024), .B1(n26132), .B2(n12930), .ZN(
        n23234) );
  OAI22_X2 U5236 ( .A1(n26325), .A2(n28025), .B1(n26131), .B2(n12930), .ZN(
        n23235) );
  OAI22_X2 U5238 ( .A1(n26325), .A2(n28026), .B1(n26279), .B2(n12930), .ZN(
        n23236) );
  OAI22_X2 U5240 ( .A1(n26325), .A2(n28027), .B1(n26278), .B2(n12930), .ZN(
        n23237) );
  OAI22_X2 U5242 ( .A1(n26325), .A2(n28028), .B1(n26277), .B2(n12930), .ZN(
        n23238) );
  OAI22_X2 U5244 ( .A1(n26325), .A2(n28029), .B1(n26276), .B2(n12930), .ZN(
        n23239) );
  OAI22_X2 U5246 ( .A1(n26325), .A2(n28030), .B1(n26275), .B2(n12930), .ZN(
        n23240) );
  OAI22_X2 U5248 ( .A1(n26325), .A2(n28031), .B1(n26274), .B2(n12930), .ZN(
        n23241) );
  OAI22_X2 U5250 ( .A1(n26325), .A2(n28032), .B1(n26273), .B2(n12930), .ZN(
        n23242) );
  OAI22_X2 U5252 ( .A1(n26325), .A2(n28033), .B1(n26272), .B2(n12930), .ZN(
        n23243) );
  OAI22_X2 U5254 ( .A1(n26325), .A2(n28034), .B1(n26271), .B2(n12930), .ZN(
        n23244) );
  OAI22_X2 U5256 ( .A1(n26325), .A2(n28035), .B1(n26270), .B2(n12930), .ZN(
        n23245) );
  OAI22_X2 U5258 ( .A1(n26325), .A2(n28036), .B1(n26269), .B2(n12930), .ZN(
        n23246) );
  OAI22_X2 U5260 ( .A1(n26325), .A2(n28037), .B1(n26268), .B2(n12930), .ZN(
        n23247) );
  OAI22_X2 U5264 ( .A1(n26324), .A2(n28038), .B1(n26134), .B2(n12948), .ZN(
        n23248) );
  OAI22_X2 U5266 ( .A1(n26324), .A2(n28039), .B1(n26133), .B2(n12948), .ZN(
        n23249) );
  OAI22_X2 U5268 ( .A1(n26324), .A2(n28040), .B1(n26132), .B2(n12948), .ZN(
        n23250) );
  OAI22_X2 U5270 ( .A1(n26324), .A2(n28041), .B1(n26131), .B2(n12948), .ZN(
        n23251) );
  OAI22_X2 U5272 ( .A1(n26324), .A2(n28042), .B1(n26279), .B2(n12948), .ZN(
        n23252) );
  OAI22_X2 U5274 ( .A1(n26324), .A2(n28043), .B1(n26278), .B2(n12948), .ZN(
        n23253) );
  OAI22_X2 U5276 ( .A1(n26324), .A2(n28044), .B1(n26277), .B2(n12948), .ZN(
        n23254) );
  OAI22_X2 U5278 ( .A1(n26324), .A2(n28045), .B1(n26276), .B2(n12948), .ZN(
        n23255) );
  OAI22_X2 U5280 ( .A1(n26324), .A2(n28046), .B1(n26275), .B2(n12948), .ZN(
        n23256) );
  OAI22_X2 U5282 ( .A1(n26324), .A2(n28047), .B1(n26274), .B2(n12948), .ZN(
        n23257) );
  OAI22_X2 U5284 ( .A1(n26324), .A2(n28048), .B1(n26273), .B2(n12948), .ZN(
        n23258) );
  OAI22_X2 U5286 ( .A1(n26324), .A2(n28049), .B1(n26272), .B2(n12948), .ZN(
        n23259) );
  OAI22_X2 U5288 ( .A1(n26324), .A2(n28050), .B1(n26271), .B2(n12948), .ZN(
        n23260) );
  OAI22_X2 U5290 ( .A1(n26324), .A2(n28051), .B1(n26270), .B2(n12948), .ZN(
        n23261) );
  OAI22_X2 U5292 ( .A1(n26324), .A2(n28052), .B1(n26269), .B2(n12948), .ZN(
        n23262) );
  OAI22_X2 U5294 ( .A1(n26324), .A2(n28053), .B1(n26268), .B2(n12948), .ZN(
        n23263) );
  NOR3_X2 U5300 ( .A1(n12967), .A2(n26502), .A3(n26506), .ZN(n12965) );
  NOR4_X2 U5302 ( .A1(n26508), .A2(n26502), .A3(n26509), .A4(n26510), .ZN(
        n12968) );
  NOR3_X2 U5304 ( .A1(n12967), .A2(n25781), .A3(n26509), .ZN(n12969) );
  NAND2_X2 U5306 ( .A1(n12971), .A2(n12972), .ZN(n12967) );
  NAND2_X2 U5310 ( .A1(n11283), .A2(n11437), .ZN(n12966) );
  OAI22_X2 U5311 ( .A1(n25958), .A2(add_1445_B_6_), .B1(n22425), .B2(n11437), 
        .ZN(n23270) );
  OAI22_X2 U5315 ( .A1(n26319), .A2(n27894), .B1(n26134), .B2(n12980), .ZN(
        n23271) );
  OAI22_X2 U5317 ( .A1(n26319), .A2(n27895), .B1(n26133), .B2(n12980), .ZN(
        n23272) );
  OAI22_X2 U5319 ( .A1(n26319), .A2(n27896), .B1(n26132), .B2(n12980), .ZN(
        n23273) );
  OAI22_X2 U5321 ( .A1(n26319), .A2(n27897), .B1(n26131), .B2(n12980), .ZN(
        n23274) );
  OAI22_X2 U5323 ( .A1(n26319), .A2(n27898), .B1(n26279), .B2(n12980), .ZN(
        n23275) );
  OAI22_X2 U5325 ( .A1(n26319), .A2(n27899), .B1(n26278), .B2(n12980), .ZN(
        n23276) );
  OAI22_X2 U5327 ( .A1(n26319), .A2(n27900), .B1(n26277), .B2(n12980), .ZN(
        n23277) );
  OAI22_X2 U5329 ( .A1(n26319), .A2(n27901), .B1(n26276), .B2(n12980), .ZN(
        n23278) );
  OAI22_X2 U5331 ( .A1(n26319), .A2(n27902), .B1(n26275), .B2(n12980), .ZN(
        n23279) );
  OAI22_X2 U5333 ( .A1(n26319), .A2(n27903), .B1(n26274), .B2(n12980), .ZN(
        n23280) );
  OAI22_X2 U5335 ( .A1(n26319), .A2(n27904), .B1(n26273), .B2(n12980), .ZN(
        n23281) );
  OAI22_X2 U5337 ( .A1(n26319), .A2(n27905), .B1(n26272), .B2(n12980), .ZN(
        n23282) );
  OAI22_X2 U5339 ( .A1(n26319), .A2(n27906), .B1(n26271), .B2(n12980), .ZN(
        n23283) );
  OAI22_X2 U5341 ( .A1(n26319), .A2(n27907), .B1(n26270), .B2(n12980), .ZN(
        n23284) );
  OAI22_X2 U5343 ( .A1(n26319), .A2(n27908), .B1(n26269), .B2(n12980), .ZN(
        n23285) );
  OAI22_X2 U5345 ( .A1(n26319), .A2(n27909), .B1(n26268), .B2(n12980), .ZN(
        n23286) );
  OAI22_X2 U5349 ( .A1(n26318), .A2(n27910), .B1(n26134), .B2(n12982), .ZN(
        n23287) );
  OAI22_X2 U5351 ( .A1(n26318), .A2(n27911), .B1(n26133), .B2(n12982), .ZN(
        n23288) );
  OAI22_X2 U5353 ( .A1(n26318), .A2(n27912), .B1(n26132), .B2(n12982), .ZN(
        n23289) );
  OAI22_X2 U5355 ( .A1(n26318), .A2(n27913), .B1(n26131), .B2(n12982), .ZN(
        n23290) );
  OAI22_X2 U5357 ( .A1(n26318), .A2(n27914), .B1(n26279), .B2(n12982), .ZN(
        n23291) );
  OAI22_X2 U5359 ( .A1(n26318), .A2(n27915), .B1(n26278), .B2(n12982), .ZN(
        n23292) );
  OAI22_X2 U5361 ( .A1(n26318), .A2(n27916), .B1(n26277), .B2(n12982), .ZN(
        n23293) );
  OAI22_X2 U5363 ( .A1(n26318), .A2(n27917), .B1(n26276), .B2(n12982), .ZN(
        n23294) );
  OAI22_X2 U5365 ( .A1(n26318), .A2(n27918), .B1(n26275), .B2(n12982), .ZN(
        n23295) );
  OAI22_X2 U5367 ( .A1(n26318), .A2(n27919), .B1(n26274), .B2(n12982), .ZN(
        n23296) );
  OAI22_X2 U5369 ( .A1(n26318), .A2(n27920), .B1(n26273), .B2(n12982), .ZN(
        n23297) );
  OAI22_X2 U5371 ( .A1(n26318), .A2(n27921), .B1(n26272), .B2(n12982), .ZN(
        n23298) );
  OAI22_X2 U5373 ( .A1(n26318), .A2(n27922), .B1(n26271), .B2(n12982), .ZN(
        n23299) );
  OAI22_X2 U5375 ( .A1(n26318), .A2(n27923), .B1(n26270), .B2(n12982), .ZN(
        n23300) );
  OAI22_X2 U5377 ( .A1(n26318), .A2(n27924), .B1(n26269), .B2(n12982), .ZN(
        n23301) );
  OAI22_X2 U5379 ( .A1(n26318), .A2(n27925), .B1(n26268), .B2(n12982), .ZN(
        n23302) );
  OAI22_X2 U5383 ( .A1(n26317), .A2(n27926), .B1(n26134), .B2(n12984), .ZN(
        n23303) );
  OAI22_X2 U5385 ( .A1(n26317), .A2(n27927), .B1(n26133), .B2(n12984), .ZN(
        n23304) );
  OAI22_X2 U5387 ( .A1(n26317), .A2(n27928), .B1(n26132), .B2(n12984), .ZN(
        n23305) );
  OAI22_X2 U5389 ( .A1(n26317), .A2(n27929), .B1(n26131), .B2(n12984), .ZN(
        n23306) );
  OAI22_X2 U5391 ( .A1(n26317), .A2(n27930), .B1(n26279), .B2(n12984), .ZN(
        n23307) );
  OAI22_X2 U5393 ( .A1(n26317), .A2(n27931), .B1(n26278), .B2(n12984), .ZN(
        n23308) );
  OAI22_X2 U5395 ( .A1(n26317), .A2(n27932), .B1(n26277), .B2(n12984), .ZN(
        n23309) );
  OAI22_X2 U5397 ( .A1(n26317), .A2(n27933), .B1(n26276), .B2(n12984), .ZN(
        n23310) );
  OAI22_X2 U5399 ( .A1(n26317), .A2(n27934), .B1(n26275), .B2(n12984), .ZN(
        n23311) );
  OAI22_X2 U5401 ( .A1(n26317), .A2(n27935), .B1(n26274), .B2(n12984), .ZN(
        n23312) );
  OAI22_X2 U5403 ( .A1(n26317), .A2(n27936), .B1(n26273), .B2(n12984), .ZN(
        n23313) );
  OAI22_X2 U5405 ( .A1(n26317), .A2(n27937), .B1(n26272), .B2(n12984), .ZN(
        n23314) );
  OAI22_X2 U5407 ( .A1(n26317), .A2(n27938), .B1(n26271), .B2(n12984), .ZN(
        n23315) );
  OAI22_X2 U5409 ( .A1(n26317), .A2(n27939), .B1(n26270), .B2(n12984), .ZN(
        n23316) );
  OAI22_X2 U5411 ( .A1(n26317), .A2(n27940), .B1(n26269), .B2(n12984), .ZN(
        n23317) );
  OAI22_X2 U5413 ( .A1(n26317), .A2(n27941), .B1(n26268), .B2(n12984), .ZN(
        n23318) );
  OAI22_X2 U5417 ( .A1(n26316), .A2(n27942), .B1(n26134), .B2(n12986), .ZN(
        n23319) );
  OAI22_X2 U5419 ( .A1(n26316), .A2(n27943), .B1(n26133), .B2(n12986), .ZN(
        n23320) );
  OAI22_X2 U5421 ( .A1(n26316), .A2(n27944), .B1(n26132), .B2(n12986), .ZN(
        n23321) );
  OAI22_X2 U5423 ( .A1(n26316), .A2(n27945), .B1(n26131), .B2(n12986), .ZN(
        n23322) );
  OAI22_X2 U5425 ( .A1(n26316), .A2(n27946), .B1(n26279), .B2(n12986), .ZN(
        n23323) );
  OAI22_X2 U5427 ( .A1(n26316), .A2(n27947), .B1(n26278), .B2(n12986), .ZN(
        n23324) );
  OAI22_X2 U5429 ( .A1(n26316), .A2(n27948), .B1(n26277), .B2(n12986), .ZN(
        n23325) );
  OAI22_X2 U5431 ( .A1(n26316), .A2(n27949), .B1(n26276), .B2(n12986), .ZN(
        n23326) );
  OAI22_X2 U5433 ( .A1(n26316), .A2(n27950), .B1(n26275), .B2(n12986), .ZN(
        n23327) );
  OAI22_X2 U5435 ( .A1(n26316), .A2(n27951), .B1(n26274), .B2(n12986), .ZN(
        n23328) );
  OAI22_X2 U5437 ( .A1(n26316), .A2(n27952), .B1(n26273), .B2(n12986), .ZN(
        n23329) );
  OAI22_X2 U5439 ( .A1(n26316), .A2(n27953), .B1(n26272), .B2(n12986), .ZN(
        n23330) );
  OAI22_X2 U5441 ( .A1(n26316), .A2(n27954), .B1(n26271), .B2(n12986), .ZN(
        n23331) );
  OAI22_X2 U5443 ( .A1(n26316), .A2(n27955), .B1(n26270), .B2(n12986), .ZN(
        n23332) );
  OAI22_X2 U5445 ( .A1(n26316), .A2(n27956), .B1(n26269), .B2(n12986), .ZN(
        n23333) );
  OAI22_X2 U5447 ( .A1(n26316), .A2(n27957), .B1(n26268), .B2(n12986), .ZN(
        n23334) );
  OAI22_X2 U5451 ( .A1(n26315), .A2(n27958), .B1(n26134), .B2(n12988), .ZN(
        n23335) );
  OAI22_X2 U5453 ( .A1(n26315), .A2(n27959), .B1(n26133), .B2(n12988), .ZN(
        n23336) );
  OAI22_X2 U5455 ( .A1(n26315), .A2(n27960), .B1(n26132), .B2(n12988), .ZN(
        n23337) );
  OAI22_X2 U5457 ( .A1(n26315), .A2(n27961), .B1(n26131), .B2(n12988), .ZN(
        n23338) );
  OAI22_X2 U5459 ( .A1(n26315), .A2(n27962), .B1(n26279), .B2(n12988), .ZN(
        n23339) );
  OAI22_X2 U5461 ( .A1(n26315), .A2(n27963), .B1(n26278), .B2(n12988), .ZN(
        n23340) );
  OAI22_X2 U5463 ( .A1(n26315), .A2(n27964), .B1(n26277), .B2(n12988), .ZN(
        n23341) );
  OAI22_X2 U5465 ( .A1(n26315), .A2(n27965), .B1(n26276), .B2(n12988), .ZN(
        n23342) );
  OAI22_X2 U5467 ( .A1(n26315), .A2(n27966), .B1(n26275), .B2(n12988), .ZN(
        n23343) );
  OAI22_X2 U5469 ( .A1(n26315), .A2(n27967), .B1(n26274), .B2(n12988), .ZN(
        n23344) );
  OAI22_X2 U5471 ( .A1(n26315), .A2(n27968), .B1(n26273), .B2(n12988), .ZN(
        n23345) );
  OAI22_X2 U5473 ( .A1(n26315), .A2(n27969), .B1(n26272), .B2(n12988), .ZN(
        n23346) );
  OAI22_X2 U5475 ( .A1(n26315), .A2(n27970), .B1(n26271), .B2(n12988), .ZN(
        n23347) );
  OAI22_X2 U5477 ( .A1(n26315), .A2(n27971), .B1(n26270), .B2(n12988), .ZN(
        n23348) );
  OAI22_X2 U5479 ( .A1(n26315), .A2(n27972), .B1(n26269), .B2(n12988), .ZN(
        n23349) );
  OAI22_X2 U5481 ( .A1(n26315), .A2(n27973), .B1(n26268), .B2(n12988), .ZN(
        n23350) );
  OAI22_X2 U5486 ( .A1(n26310), .A2(n27814), .B1(n26134), .B2(n12992), .ZN(
        n23351) );
  OAI22_X2 U5488 ( .A1(n26310), .A2(n27815), .B1(n26133), .B2(n12992), .ZN(
        n23352) );
  OAI22_X2 U5490 ( .A1(n26310), .A2(n27816), .B1(n26132), .B2(n12992), .ZN(
        n23353) );
  OAI22_X2 U5492 ( .A1(n26310), .A2(n27817), .B1(n26131), .B2(n12992), .ZN(
        n23354) );
  OAI22_X2 U5494 ( .A1(n26310), .A2(n27818), .B1(n26279), .B2(n12992), .ZN(
        n23355) );
  OAI22_X2 U5496 ( .A1(n26310), .A2(n27819), .B1(n26278), .B2(n12992), .ZN(
        n23356) );
  OAI22_X2 U5498 ( .A1(n26310), .A2(n27820), .B1(n26277), .B2(n12992), .ZN(
        n23357) );
  OAI22_X2 U5500 ( .A1(n26310), .A2(n27821), .B1(n26276), .B2(n12992), .ZN(
        n23358) );
  OAI22_X2 U5502 ( .A1(n26310), .A2(n27822), .B1(n26275), .B2(n12992), .ZN(
        n23359) );
  OAI22_X2 U5504 ( .A1(n26310), .A2(n27823), .B1(n26274), .B2(n12992), .ZN(
        n23360) );
  OAI22_X2 U5506 ( .A1(n26310), .A2(n27824), .B1(n26273), .B2(n12992), .ZN(
        n23361) );
  OAI22_X2 U5508 ( .A1(n26310), .A2(n27825), .B1(n26272), .B2(n12992), .ZN(
        n23362) );
  OAI22_X2 U5510 ( .A1(n26310), .A2(n27826), .B1(n26271), .B2(n12992), .ZN(
        n23363) );
  OAI22_X2 U5512 ( .A1(n26310), .A2(n27827), .B1(n26270), .B2(n12992), .ZN(
        n23364) );
  OAI22_X2 U5514 ( .A1(n26310), .A2(n27828), .B1(n26269), .B2(n12992), .ZN(
        n23365) );
  OAI22_X2 U5516 ( .A1(n26310), .A2(n27829), .B1(n26268), .B2(n12992), .ZN(
        n23366) );
  OAI22_X2 U5520 ( .A1(n26309), .A2(n27830), .B1(n26134), .B2(n13009), .ZN(
        n23367) );
  OAI22_X2 U5522 ( .A1(n26309), .A2(n27831), .B1(n26133), .B2(n13009), .ZN(
        n23368) );
  OAI22_X2 U5524 ( .A1(n26309), .A2(n27832), .B1(n26132), .B2(n13009), .ZN(
        n23369) );
  OAI22_X2 U5526 ( .A1(n26309), .A2(n27833), .B1(n26131), .B2(n13009), .ZN(
        n23370) );
  OAI22_X2 U5528 ( .A1(n26309), .A2(n27834), .B1(n26279), .B2(n13009), .ZN(
        n23371) );
  OAI22_X2 U5530 ( .A1(n26309), .A2(n27835), .B1(n26278), .B2(n13009), .ZN(
        n23372) );
  OAI22_X2 U5532 ( .A1(n26309), .A2(n27836), .B1(n26277), .B2(n13009), .ZN(
        n23373) );
  OAI22_X2 U5534 ( .A1(n26309), .A2(n27837), .B1(n26276), .B2(n13009), .ZN(
        n23374) );
  OAI22_X2 U5536 ( .A1(n26309), .A2(n27838), .B1(n26275), .B2(n13009), .ZN(
        n23375) );
  OAI22_X2 U5538 ( .A1(n26309), .A2(n27839), .B1(n26274), .B2(n13009), .ZN(
        n23376) );
  OAI22_X2 U5540 ( .A1(n26309), .A2(n27840), .B1(n26273), .B2(n13009), .ZN(
        n23377) );
  OAI22_X2 U5542 ( .A1(n26309), .A2(n27841), .B1(n26272), .B2(n13009), .ZN(
        n23378) );
  OAI22_X2 U5544 ( .A1(n26309), .A2(n27842), .B1(n26271), .B2(n13009), .ZN(
        n23379) );
  OAI22_X2 U5546 ( .A1(n26309), .A2(n27843), .B1(n26270), .B2(n13009), .ZN(
        n23380) );
  OAI22_X2 U5548 ( .A1(n26309), .A2(n27844), .B1(n26269), .B2(n13009), .ZN(
        n23381) );
  OAI22_X2 U5550 ( .A1(n26309), .A2(n27845), .B1(n26268), .B2(n13009), .ZN(
        n23382) );
  OAI22_X2 U5554 ( .A1(n26308), .A2(n27846), .B1(n26134), .B2(n13012), .ZN(
        n23383) );
  OAI22_X2 U5556 ( .A1(n26308), .A2(n27847), .B1(n26133), .B2(n13012), .ZN(
        n23384) );
  OAI22_X2 U5558 ( .A1(n26308), .A2(n27848), .B1(n26132), .B2(n13012), .ZN(
        n23385) );
  OAI22_X2 U5560 ( .A1(n26308), .A2(n27849), .B1(n26131), .B2(n13012), .ZN(
        n23386) );
  OAI22_X2 U5562 ( .A1(n26308), .A2(n27850), .B1(n26279), .B2(n13012), .ZN(
        n23387) );
  OAI22_X2 U5564 ( .A1(n26308), .A2(n27851), .B1(n26278), .B2(n13012), .ZN(
        n23388) );
  OAI22_X2 U5566 ( .A1(n26308), .A2(n27852), .B1(n26277), .B2(n13012), .ZN(
        n23389) );
  OAI22_X2 U5568 ( .A1(n26308), .A2(n27853), .B1(n26276), .B2(n13012), .ZN(
        n23390) );
  OAI22_X2 U5570 ( .A1(n26308), .A2(n27854), .B1(n26275), .B2(n13012), .ZN(
        n23391) );
  OAI22_X2 U5572 ( .A1(n26308), .A2(n27855), .B1(n26274), .B2(n13012), .ZN(
        n23392) );
  OAI22_X2 U5574 ( .A1(n26308), .A2(n27856), .B1(n26273), .B2(n13012), .ZN(
        n23393) );
  OAI22_X2 U5576 ( .A1(n26308), .A2(n27857), .B1(n26272), .B2(n13012), .ZN(
        n23394) );
  OAI22_X2 U5578 ( .A1(n26308), .A2(n27858), .B1(n26271), .B2(n13012), .ZN(
        n23395) );
  OAI22_X2 U5580 ( .A1(n26308), .A2(n27859), .B1(n26270), .B2(n13012), .ZN(
        n23396) );
  OAI22_X2 U5582 ( .A1(n26308), .A2(n27860), .B1(n26269), .B2(n13012), .ZN(
        n23397) );
  OAI22_X2 U5584 ( .A1(n26308), .A2(n27861), .B1(n26268), .B2(n13012), .ZN(
        n23398) );
  OAI22_X2 U5588 ( .A1(n26307), .A2(n27862), .B1(n26134), .B2(n13029), .ZN(
        n23399) );
  OAI22_X2 U5590 ( .A1(n26307), .A2(n27863), .B1(n26133), .B2(n13029), .ZN(
        n23400) );
  OAI22_X2 U5592 ( .A1(n26307), .A2(n27864), .B1(n26132), .B2(n13029), .ZN(
        n23401) );
  OAI22_X2 U5594 ( .A1(n26307), .A2(n27865), .B1(n26131), .B2(n13029), .ZN(
        n23402) );
  OAI22_X2 U5596 ( .A1(n26307), .A2(n27866), .B1(n26279), .B2(n13029), .ZN(
        n23403) );
  OAI22_X2 U5598 ( .A1(n26307), .A2(n27867), .B1(n26278), .B2(n13029), .ZN(
        n23404) );
  OAI22_X2 U5600 ( .A1(n26307), .A2(n27868), .B1(n26277), .B2(n13029), .ZN(
        n23405) );
  OAI22_X2 U5602 ( .A1(n26307), .A2(n27869), .B1(n26276), .B2(n13029), .ZN(
        n23406) );
  OAI22_X2 U5604 ( .A1(n26307), .A2(n27870), .B1(n26275), .B2(n13029), .ZN(
        n23407) );
  OAI22_X2 U5606 ( .A1(n26307), .A2(n27871), .B1(n26274), .B2(n13029), .ZN(
        n23408) );
  OAI22_X2 U5608 ( .A1(n26307), .A2(n27872), .B1(n26273), .B2(n13029), .ZN(
        n23409) );
  OAI22_X2 U5610 ( .A1(n26307), .A2(n27873), .B1(n26272), .B2(n13029), .ZN(
        n23410) );
  OAI22_X2 U5612 ( .A1(n26307), .A2(n27874), .B1(n26271), .B2(n13029), .ZN(
        n23411) );
  OAI22_X2 U5614 ( .A1(n26307), .A2(n27875), .B1(n26270), .B2(n13029), .ZN(
        n23412) );
  OAI22_X2 U5616 ( .A1(n26307), .A2(n27876), .B1(n26269), .B2(n13029), .ZN(
        n23413) );
  OAI22_X2 U5618 ( .A1(n26307), .A2(n27877), .B1(n26268), .B2(n13029), .ZN(
        n23414) );
  OAI22_X2 U5622 ( .A1(n26306), .A2(n27878), .B1(n26134), .B2(n13031), .ZN(
        n23415) );
  OAI22_X2 U5625 ( .A1(n26306), .A2(n27879), .B1(n26133), .B2(n13031), .ZN(
        n23416) );
  OAI22_X2 U5628 ( .A1(n26306), .A2(n27880), .B1(n26132), .B2(n13031), .ZN(
        n23417) );
  OAI22_X2 U5631 ( .A1(n26306), .A2(n27881), .B1(n26131), .B2(n13031), .ZN(
        n23418) );
  OAI22_X2 U5634 ( .A1(n26306), .A2(n27882), .B1(n26279), .B2(n13031), .ZN(
        n23419) );
  OAI22_X2 U5637 ( .A1(n26306), .A2(n27883), .B1(n26278), .B2(n13031), .ZN(
        n23420) );
  OAI22_X2 U5640 ( .A1(n26306), .A2(n27884), .B1(n26277), .B2(n13031), .ZN(
        n23421) );
  OAI22_X2 U5643 ( .A1(n26306), .A2(n27885), .B1(n26276), .B2(n13031), .ZN(
        n23422) );
  OAI22_X2 U5646 ( .A1(n26306), .A2(n27886), .B1(n26275), .B2(n13031), .ZN(
        n23423) );
  OAI22_X2 U5649 ( .A1(n26306), .A2(n27887), .B1(n26274), .B2(n13031), .ZN(
        n23424) );
  OAI22_X2 U5652 ( .A1(n26306), .A2(n27888), .B1(n26273), .B2(n13031), .ZN(
        n23425) );
  OAI22_X2 U5655 ( .A1(n26306), .A2(n27889), .B1(n26272), .B2(n13031), .ZN(
        n23426) );
  OAI22_X2 U5658 ( .A1(n26306), .A2(n27890), .B1(n26271), .B2(n13031), .ZN(
        n23427) );
  OAI22_X2 U5661 ( .A1(n26306), .A2(n27891), .B1(n26270), .B2(n13031), .ZN(
        n23428) );
  OAI22_X2 U5664 ( .A1(n26306), .A2(n27892), .B1(n26269), .B2(n13031), .ZN(
        n23429) );
  OAI22_X2 U5667 ( .A1(n26306), .A2(n27893), .B1(n26268), .B2(n13031), .ZN(
        n23430) );
  AND3_X2 U5673 ( .A1(n22426), .A2(n26135), .A3(n16374), .ZN(n11794) );
  NAND2_X2 U5688 ( .A1(n13045), .A2(n13046), .ZN(n23434) );
  NAND3_X2 U5689 ( .A1(n26302), .A2(n22414), .A3(add_283_carry[5]), .ZN(n13046) );
  OAI22_X2 U5708 ( .A1(n22419), .A2(n13054), .B1(add_283_A_0_), .B2(n13055), 
        .ZN(n23439) );
  NAND3_X2 U5709 ( .A1(n13054), .A2(n11878), .A3(n11634), .ZN(n13055) );
  NAND2_X2 U5711 ( .A1(n11634), .A2(n10081), .ZN(n13054) );
  NAND2_X2 U5716 ( .A1(n13057), .A2(n13058), .ZN(n23441) );
  NAND3_X2 U5717 ( .A1(add_262_carry[9]), .A2(n13059), .A3(n22407), .ZN(n13058) );
  NOR3_X2 U5719 ( .A1(n26293), .A2(add_262_carry[9]), .A3(n13063), .ZN(n13060)
         );
  OAI22_X2 U5720 ( .A1(n22413), .A2(n11441), .B1(add_1445_B_0_), .B2(n26280), 
        .ZN(n23442) );
  NOR3_X2 U5722 ( .A1(n13063), .A2(n26296), .A3(n26293), .ZN(n13059) );
  AND4_X2 U5724 ( .A1(n22410), .A2(n22411), .A3(n13065), .A4(n13066), .ZN(
        n13063) );
  AND3_X2 U5725 ( .A1(n13067), .A2(n18745), .A3(n18744), .ZN(n13066) );
  AND3_X2 U5726 ( .A1(n22408), .A2(n22409), .A3(n25775), .ZN(n13067) );
  AND3_X2 U5727 ( .A1(n22412), .A2(add_1445_B_9_), .A3(n22413), .ZN(n13065) );
  NOR2_X2 U5731 ( .A1(n13068), .A2(n26293), .ZN(n23443) );
  AND3_X2 U5735 ( .A1(n24896), .A2(n25257), .A3(n12146), .ZN(n12057) );
  NOR3_X2 U5736 ( .A1(n26350), .A2(n22399), .A3(n26137), .ZN(n12146) );
  OAI22_X2 U5737 ( .A1(n22400), .A2(n26293), .B1(n11399), .B2(n13071), .ZN(
        n23444) );
  NAND4_X2 U5742 ( .A1(n26138), .A2(n11634), .A3(n13075), .A4(n25253), .ZN(
        n11399) );
  NAND2_X2 U5750 ( .A1(n13069), .A2(n13080), .ZN(n13078) );
  NAND3_X2 U5751 ( .A1(n24896), .A2(n25257), .A3(n24865), .ZN(n13080) );
  OAI22_X2 U5759 ( .A1(n22404), .A2(n26282), .B1(n13084), .B2(n13088), .ZN(
        n23448) );
  OAI22_X2 U5763 ( .A1(n22405), .A2(n13091), .B1(n25104), .B2(n13084), .ZN(
        n23449) );
  OAI22_X2 U5768 ( .A1(n22406), .A2(n13075), .B1(n26283), .B2(n13092), .ZN(
        n23450) );
  NOR2_X2 U5771 ( .A1(n26293), .A2(n13069), .ZN(n13085) );
  AND4_X2 U5772 ( .A1(n18743), .A2(n22404), .A3(n22405), .A4(n22406), .ZN(
        n13069) );
  OAI22_X2 U5775 ( .A1(n26294), .A2(n26293), .B1(n22399), .B2(n13095), .ZN(
        n23451) );
  NAND2_X2 U5777 ( .A1(n11634), .A2(n13096), .ZN(n13095) );
  NAND3_X2 U5778 ( .A1(n12803), .A2(n26135), .A3(n27801), .ZN(n13096) );
  NAND4_X2 U5782 ( .A1(n13101), .A2(n13102), .A3(n13103), .A4(n13104), .ZN(
        n13100) );
  AOI221_X2 U5783 ( .B1(n25905), .B2(n25052), .C1(n25904), .C2(n25551), .A(
        n13109), .ZN(n13104) );
  AOI221_X2 U5787 ( .B1(n25895), .B2(n25051), .C1(n25894), .C2(n25550), .A(
        n13119), .ZN(n13103) );
  OAI22_X2 U5788 ( .A1(n18736), .A2(n25891), .B1(n18708), .B2(n25889), .ZN(
        n13119) );
  AOI221_X2 U5791 ( .B1(n18721), .B2(n25888), .C1(n18712), .C2(n25885), .A(
        n13124), .ZN(n13102) );
  AOI221_X2 U5793 ( .B1(n18738), .B2(n25877), .C1(n18729), .C2(n25876), .A(
        n13132), .ZN(n13101) );
  OAI22_X2 U5794 ( .A1(n25873), .A2(n26663), .B1(n25871), .B2(n26679), .ZN(
        n13132) );
  NAND4_X2 U5795 ( .A1(n13137), .A2(n13138), .A3(n13139), .A4(n13140), .ZN(
        n13099) );
  AOI221_X2 U5796 ( .B1(n18710), .B2(n25869), .C1(n25868), .C2(n25549), .A(
        n13144), .ZN(n13140) );
  AOI221_X2 U5799 ( .B1(n25859), .B2(n25697), .C1(n25858), .C2(n25210), .A(
        n13155), .ZN(n13139) );
  OAI22_X2 U5800 ( .A1(n18741), .A2(n25855), .B1(n18713), .B2(n25853), .ZN(
        n13155) );
  AOI221_X2 U5803 ( .B1(n18733), .B2(n25851), .C1(n18724), .C2(n25850), .A(
        n13160), .ZN(n13138) );
  AOI221_X2 U5805 ( .B1(n18734), .B2(n25841), .C1(n18725), .C2(n25840), .A(
        n13166), .ZN(n13137) );
  OAI22_X2 U5806 ( .A1(n25837), .A2(n27127), .B1(n25835), .B2(n27191), .ZN(
        n13166) );
  NAND4_X2 U5809 ( .A1(n13174), .A2(n13175), .A3(n13176), .A4(n13177), .ZN(
        n13173) );
  AOI221_X2 U5810 ( .B1(n25905), .B2(n25050), .C1(n25903), .C2(n25548), .A(
        n13180), .ZN(n13177) );
  AOI221_X2 U5814 ( .B1(n25895), .B2(n25049), .C1(n25893), .C2(n25547), .A(
        n13185), .ZN(n13176) );
  OAI22_X2 U5815 ( .A1(n18699), .A2(n25891), .B1(n18671), .B2(n25889), .ZN(
        n13185) );
  AOI221_X2 U5818 ( .B1(n18684), .B2(n25887), .C1(n18675), .C2(n25886), .A(
        n13186), .ZN(n13175) );
  AOI221_X2 U5820 ( .B1(n18701), .B2(n25877), .C1(n18692), .C2(n25875), .A(
        n13189), .ZN(n13174) );
  OAI22_X2 U5821 ( .A1(n25873), .A2(n26664), .B1(n25872), .B2(n26680), .ZN(
        n13189) );
  NAND4_X2 U5822 ( .A1(n13192), .A2(n13193), .A3(n13194), .A4(n13195), .ZN(
        n13172) );
  AOI221_X2 U5823 ( .B1(n18673), .B2(n25870), .C1(n25867), .C2(n25546), .A(
        n13197), .ZN(n13195) );
  AOI221_X2 U5826 ( .B1(n25859), .B2(n25696), .C1(n25857), .C2(n25209), .A(
        n13203), .ZN(n13194) );
  OAI22_X2 U5827 ( .A1(n18704), .A2(n25855), .B1(n18676), .B2(n25853), .ZN(
        n13203) );
  AOI221_X2 U5830 ( .B1(n18696), .B2(n25851), .C1(n18687), .C2(n25849), .A(
        n13204), .ZN(n13193) );
  AOI221_X2 U5832 ( .B1(n18697), .B2(n25841), .C1(n18688), .C2(n25839), .A(
        n13205), .ZN(n13192) );
  OAI22_X2 U5833 ( .A1(n25837), .A2(n27128), .B1(n25835), .B2(n27192), .ZN(
        n13205) );
  NAND4_X2 U5836 ( .A1(n13211), .A2(n13212), .A3(n13213), .A4(n13214), .ZN(
        n13210) );
  AOI221_X2 U5837 ( .B1(n25905), .B2(n25048), .C1(n25904), .C2(n25545), .A(
        n13217), .ZN(n13214) );
  AOI221_X2 U5841 ( .B1(n25895), .B2(n25047), .C1(n25894), .C2(n25544), .A(
        n13222), .ZN(n13213) );
  OAI22_X2 U5842 ( .A1(n18662), .A2(n25891), .B1(n18634), .B2(n25890), .ZN(
        n13222) );
  AOI221_X2 U5845 ( .B1(n18647), .B2(n25888), .C1(n18638), .C2(n25886), .A(
        n13223), .ZN(n13212) );
  AOI221_X2 U5847 ( .B1(n18664), .B2(n25877), .C1(n18655), .C2(n25876), .A(
        n13226), .ZN(n13211) );
  OAI22_X2 U5848 ( .A1(n25873), .A2(n26665), .B1(n25871), .B2(n26681), .ZN(
        n13226) );
  NAND4_X2 U5849 ( .A1(n13229), .A2(n13230), .A3(n13231), .A4(n13232), .ZN(
        n13209) );
  AOI221_X2 U5850 ( .B1(n18636), .B2(n25869), .C1(n25868), .C2(n25543), .A(
        n13234), .ZN(n13232) );
  AOI221_X2 U5853 ( .B1(n25859), .B2(n25695), .C1(n25858), .C2(n25208), .A(
        n13240), .ZN(n13231) );
  OAI22_X2 U5854 ( .A1(n18667), .A2(n25855), .B1(n18639), .B2(n25854), .ZN(
        n13240) );
  AOI221_X2 U5857 ( .B1(n18659), .B2(n25851), .C1(n18650), .C2(n25850), .A(
        n13241), .ZN(n13230) );
  AOI221_X2 U5859 ( .B1(n18660), .B2(n25841), .C1(n18651), .C2(n25840), .A(
        n13242), .ZN(n13229) );
  OAI22_X2 U5860 ( .A1(n25837), .A2(n27129), .B1(n25835), .B2(n27193), .ZN(
        n13242) );
  NAND4_X2 U5863 ( .A1(n13248), .A2(n13249), .A3(n13250), .A4(n13251), .ZN(
        n13247) );
  AOI221_X2 U5864 ( .B1(n25905), .B2(n25046), .C1(n25903), .C2(n25542), .A(
        n13254), .ZN(n13251) );
  AOI221_X2 U5868 ( .B1(n25895), .B2(n25045), .C1(n25893), .C2(n25541), .A(
        n13259), .ZN(n13250) );
  OAI22_X2 U5869 ( .A1(n18625), .A2(n25891), .B1(n18597), .B2(n25889), .ZN(
        n13259) );
  AOI221_X2 U5872 ( .B1(n18610), .B2(n25887), .C1(n18601), .C2(n25886), .A(
        n13260), .ZN(n13249) );
  AOI221_X2 U5874 ( .B1(n18627), .B2(n25877), .C1(n18618), .C2(n25875), .A(
        n13263), .ZN(n13248) );
  OAI22_X2 U5875 ( .A1(n25873), .A2(n26666), .B1(n25871), .B2(n26682), .ZN(
        n13263) );
  NAND4_X2 U5876 ( .A1(n13266), .A2(n13267), .A3(n13268), .A4(n13269), .ZN(
        n13246) );
  AOI221_X2 U5877 ( .B1(n18599), .B2(n25870), .C1(n25868), .C2(n25540), .A(
        n13271), .ZN(n13269) );
  AOI221_X2 U5880 ( .B1(n25859), .B2(n25694), .C1(n25857), .C2(n25207), .A(
        n13277), .ZN(n13268) );
  OAI22_X2 U5881 ( .A1(n18630), .A2(n25855), .B1(n18602), .B2(n25853), .ZN(
        n13277) );
  AOI221_X2 U5884 ( .B1(n18622), .B2(n25851), .C1(n18613), .C2(n25850), .A(
        n13278), .ZN(n13267) );
  AOI221_X2 U5886 ( .B1(n18623), .B2(n25841), .C1(n18614), .C2(n25839), .A(
        n13279), .ZN(n13266) );
  OAI22_X2 U5887 ( .A1(n25837), .A2(n27130), .B1(n25836), .B2(n27194), .ZN(
        n13279) );
  NAND4_X2 U5890 ( .A1(n13285), .A2(n13286), .A3(n13287), .A4(n13288), .ZN(
        n13284) );
  AOI221_X2 U5891 ( .B1(n25905), .B2(n25044), .C1(n25904), .C2(n25539), .A(
        n13291), .ZN(n13288) );
  AOI221_X2 U5895 ( .B1(n25895), .B2(n25043), .C1(n25893), .C2(n25538), .A(
        n13296), .ZN(n13287) );
  OAI22_X2 U5896 ( .A1(n18588), .A2(n25891), .B1(n18560), .B2(n25889), .ZN(
        n13296) );
  AOI221_X2 U5899 ( .B1(n18573), .B2(n25888), .C1(n18564), .C2(n25885), .A(
        n13297), .ZN(n13286) );
  AOI221_X2 U5901 ( .B1(n18590), .B2(n25877), .C1(n18581), .C2(n25876), .A(
        n13300), .ZN(n13285) );
  OAI22_X2 U5902 ( .A1(n25873), .A2(n26667), .B1(n25871), .B2(n26683), .ZN(
        n13300) );
  NAND4_X2 U5903 ( .A1(n13303), .A2(n13304), .A3(n13305), .A4(n13306), .ZN(
        n13283) );
  AOI221_X2 U5904 ( .B1(n18562), .B2(n25869), .C1(n25867), .C2(n25537), .A(
        n13308), .ZN(n13306) );
  AOI221_X2 U5907 ( .B1(n25859), .B2(n25693), .C1(n25858), .C2(n25206), .A(
        n13314), .ZN(n13305) );
  OAI22_X2 U5908 ( .A1(n18593), .A2(n25855), .B1(n18565), .B2(n25853), .ZN(
        n13314) );
  AOI221_X2 U5911 ( .B1(n18585), .B2(n25851), .C1(n18576), .C2(n25849), .A(
        n13315), .ZN(n13304) );
  AOI221_X2 U5913 ( .B1(n18586), .B2(n25841), .C1(n18577), .C2(n25840), .A(
        n13316), .ZN(n13303) );
  OAI22_X2 U5914 ( .A1(n25837), .A2(n27131), .B1(n25835), .B2(n27195), .ZN(
        n13316) );
  NAND4_X2 U5917 ( .A1(n13322), .A2(n13323), .A3(n13324), .A4(n13325), .ZN(
        n13321) );
  AOI221_X2 U5918 ( .B1(n25905), .B2(n25042), .C1(n25903), .C2(n25536), .A(
        n13328), .ZN(n13325) );
  AOI221_X2 U5922 ( .B1(n25895), .B2(n25041), .C1(n25893), .C2(n25535), .A(
        n13333), .ZN(n13324) );
  OAI22_X2 U5923 ( .A1(n18551), .A2(n25891), .B1(n18523), .B2(n25889), .ZN(
        n13333) );
  AOI221_X2 U5926 ( .B1(n18536), .B2(n25887), .C1(n18527), .C2(n25886), .A(
        n13334), .ZN(n13323) );
  AOI221_X2 U5928 ( .B1(n18553), .B2(n25877), .C1(n18544), .C2(n25875), .A(
        n13337), .ZN(n13322) );
  OAI22_X2 U5929 ( .A1(n25873), .A2(n26668), .B1(n25872), .B2(n26684), .ZN(
        n13337) );
  NAND4_X2 U5930 ( .A1(n13340), .A2(n13341), .A3(n13342), .A4(n13343), .ZN(
        n13320) );
  AOI221_X2 U5931 ( .B1(n18525), .B2(n25870), .C1(n25867), .C2(n25534), .A(
        n13345), .ZN(n13343) );
  AOI221_X2 U5934 ( .B1(n25859), .B2(n25692), .C1(n25857), .C2(n25205), .A(
        n13351), .ZN(n13342) );
  OAI22_X2 U5935 ( .A1(n18556), .A2(n25855), .B1(n18528), .B2(n25853), .ZN(
        n13351) );
  AOI221_X2 U5938 ( .B1(n18548), .B2(n25851), .C1(n18539), .C2(n25849), .A(
        n13352), .ZN(n13341) );
  AOI221_X2 U5940 ( .B1(n18549), .B2(n25841), .C1(n18540), .C2(n25839), .A(
        n13353), .ZN(n13340) );
  OAI22_X2 U5941 ( .A1(n25837), .A2(n27132), .B1(n25835), .B2(n27196), .ZN(
        n13353) );
  NAND4_X2 U5944 ( .A1(n13359), .A2(n13360), .A3(n13361), .A4(n13362), .ZN(
        n13358) );
  AOI221_X2 U5945 ( .B1(n25905), .B2(n25040), .C1(n25904), .C2(n25533), .A(
        n13365), .ZN(n13362) );
  AOI221_X2 U5949 ( .B1(n25895), .B2(n25039), .C1(n25894), .C2(n25532), .A(
        n13370), .ZN(n13361) );
  OAI22_X2 U5950 ( .A1(n18514), .A2(n25891), .B1(n18486), .B2(n25890), .ZN(
        n13370) );
  AOI221_X2 U5953 ( .B1(n18499), .B2(n25888), .C1(n18490), .C2(n25885), .A(
        n13371), .ZN(n13360) );
  AOI221_X2 U5955 ( .B1(n18516), .B2(n25877), .C1(n18507), .C2(n25876), .A(
        n13374), .ZN(n13359) );
  OAI22_X2 U5956 ( .A1(n25873), .A2(n26669), .B1(n25871), .B2(n26685), .ZN(
        n13374) );
  NAND4_X2 U5957 ( .A1(n13377), .A2(n13378), .A3(n13379), .A4(n13380), .ZN(
        n13357) );
  AOI221_X2 U5958 ( .B1(n18488), .B2(n25869), .C1(n25868), .C2(n25531), .A(
        n13382), .ZN(n13380) );
  AOI221_X2 U5961 ( .B1(n25859), .B2(n25691), .C1(n25858), .C2(n25204), .A(
        n13388), .ZN(n13379) );
  OAI22_X2 U5962 ( .A1(n18519), .A2(n25855), .B1(n18491), .B2(n25854), .ZN(
        n13388) );
  AOI221_X2 U5965 ( .B1(n18511), .B2(n25851), .C1(n18502), .C2(n25850), .A(
        n13389), .ZN(n13378) );
  AOI221_X2 U5967 ( .B1(n18512), .B2(n25841), .C1(n18503), .C2(n25840), .A(
        n13390), .ZN(n13377) );
  OAI22_X2 U5968 ( .A1(n25837), .A2(n27133), .B1(n25835), .B2(n27197), .ZN(
        n13390) );
  NAND4_X2 U5971 ( .A1(n13396), .A2(n13397), .A3(n13398), .A4(n13399), .ZN(
        n13395) );
  AOI221_X2 U5972 ( .B1(n25905), .B2(n25038), .C1(n25904), .C2(n25530), .A(
        n13402), .ZN(n13399) );
  AOI221_X2 U5976 ( .B1(n25895), .B2(n25037), .C1(n25894), .C2(n25529), .A(
        n13407), .ZN(n13398) );
  OAI22_X2 U5977 ( .A1(n18477), .A2(n25891), .B1(n18449), .B2(n25889), .ZN(
        n13407) );
  AOI221_X2 U5980 ( .B1(n18462), .B2(n25888), .C1(n18453), .C2(n25886), .A(
        n13408), .ZN(n13397) );
  AOI221_X2 U5982 ( .B1(n18479), .B2(n25877), .C1(n18470), .C2(n25876), .A(
        n13411), .ZN(n13396) );
  OAI22_X2 U5983 ( .A1(n25873), .A2(n26670), .B1(n25872), .B2(n26686), .ZN(
        n13411) );
  NAND4_X2 U5984 ( .A1(n13414), .A2(n13415), .A3(n13416), .A4(n13417), .ZN(
        n13394) );
  AOI221_X2 U5985 ( .B1(n18451), .B2(n25870), .C1(n25868), .C2(n25528), .A(
        n13419), .ZN(n13417) );
  AOI221_X2 U5988 ( .B1(n25859), .B2(n25690), .C1(n25858), .C2(n25203), .A(
        n13425), .ZN(n13416) );
  OAI22_X2 U5989 ( .A1(n18482), .A2(n25855), .B1(n18454), .B2(n25853), .ZN(
        n13425) );
  AOI221_X2 U5992 ( .B1(n18474), .B2(n25851), .C1(n18465), .C2(n25850), .A(
        n13426), .ZN(n13415) );
  AOI221_X2 U5994 ( .B1(n18475), .B2(n25841), .C1(n18466), .C2(n25840), .A(
        n13427), .ZN(n13414) );
  OAI22_X2 U5995 ( .A1(n25837), .A2(n27134), .B1(n25835), .B2(n27198), .ZN(
        n13427) );
  NAND4_X2 U5998 ( .A1(n13433), .A2(n13434), .A3(n13435), .A4(n13436), .ZN(
        n13432) );
  AOI221_X2 U5999 ( .B1(n25905), .B2(n25036), .C1(n25904), .C2(n25527), .A(
        n13439), .ZN(n13436) );
  AOI221_X2 U6003 ( .B1(n25895), .B2(n25035), .C1(n25894), .C2(n25526), .A(
        n13444), .ZN(n13435) );
  OAI22_X2 U6004 ( .A1(n18440), .A2(n25891), .B1(n18412), .B2(n25889), .ZN(
        n13444) );
  AOI221_X2 U6007 ( .B1(n18425), .B2(n25887), .C1(n18416), .C2(n25885), .A(
        n13445), .ZN(n13434) );
  AOI221_X2 U6009 ( .B1(n18442), .B2(n25877), .C1(n18433), .C2(n25876), .A(
        n13448), .ZN(n13433) );
  OAI22_X2 U6010 ( .A1(n25873), .A2(n26671), .B1(n25871), .B2(n26687), .ZN(
        n13448) );
  NAND4_X2 U6011 ( .A1(n13451), .A2(n13452), .A3(n13453), .A4(n13454), .ZN(
        n13431) );
  AOI221_X2 U6012 ( .B1(n18414), .B2(n25869), .C1(n25868), .C2(n25525), .A(
        n13456), .ZN(n13454) );
  AOI221_X2 U6015 ( .B1(n25859), .B2(n25689), .C1(n25858), .C2(n25202), .A(
        n13462), .ZN(n13453) );
  OAI22_X2 U6016 ( .A1(n18445), .A2(n25855), .B1(n18417), .B2(n25853), .ZN(
        n13462) );
  AOI221_X2 U6019 ( .B1(n18437), .B2(n25851), .C1(n18428), .C2(n25850), .A(
        n13463), .ZN(n13452) );
  AOI221_X2 U6021 ( .B1(n18438), .B2(n25841), .C1(n18429), .C2(n25840), .A(
        n13464), .ZN(n13451) );
  OAI22_X2 U6022 ( .A1(n25837), .A2(n27135), .B1(n25835), .B2(n27199), .ZN(
        n13464) );
  NAND4_X2 U6025 ( .A1(n13470), .A2(n13471), .A3(n13472), .A4(n13473), .ZN(
        n13469) );
  AOI221_X2 U6026 ( .B1(n25905), .B2(n25034), .C1(n25903), .C2(n25524), .A(
        n13476), .ZN(n13473) );
  AOI221_X2 U6030 ( .B1(n25895), .B2(n25033), .C1(n25893), .C2(n25523), .A(
        n13481), .ZN(n13472) );
  OAI22_X2 U6031 ( .A1(n18403), .A2(n25891), .B1(n18375), .B2(n25889), .ZN(
        n13481) );
  AOI221_X2 U6034 ( .B1(n18388), .B2(n25888), .C1(n18379), .C2(n25886), .A(
        n13482), .ZN(n13471) );
  AOI221_X2 U6036 ( .B1(n18405), .B2(n25877), .C1(n18396), .C2(n25875), .A(
        n13485), .ZN(n13470) );
  OAI22_X2 U6037 ( .A1(n25873), .A2(n26672), .B1(n25871), .B2(n26688), .ZN(
        n13485) );
  NAND4_X2 U6038 ( .A1(n13488), .A2(n13489), .A3(n13490), .A4(n13491), .ZN(
        n13468) );
  AOI221_X2 U6039 ( .B1(n18377), .B2(n25870), .C1(n25867), .C2(n25522), .A(
        n13493), .ZN(n13491) );
  AOI221_X2 U6042 ( .B1(n25859), .B2(n25688), .C1(n25857), .C2(n25201), .A(
        n13499), .ZN(n13490) );
  OAI22_X2 U6043 ( .A1(n18408), .A2(n25855), .B1(n18380), .B2(n25853), .ZN(
        n13499) );
  AOI221_X2 U6046 ( .B1(n18400), .B2(n25851), .C1(n18391), .C2(n25849), .A(
        n13500), .ZN(n13489) );
  AOI221_X2 U6048 ( .B1(n18401), .B2(n25841), .C1(n18392), .C2(n25839), .A(
        n13501), .ZN(n13488) );
  OAI22_X2 U6049 ( .A1(n25837), .A2(n27136), .B1(n25836), .B2(n27200), .ZN(
        n13501) );
  NAND4_X2 U6052 ( .A1(n13507), .A2(n13508), .A3(n13509), .A4(n13510), .ZN(
        n13506) );
  AOI221_X2 U6053 ( .B1(n25905), .B2(n25032), .C1(n25904), .C2(n25521), .A(
        n13513), .ZN(n13510) );
  AOI221_X2 U6057 ( .B1(n25895), .B2(n25031), .C1(n25894), .C2(n25520), .A(
        n13518), .ZN(n13509) );
  OAI22_X2 U6058 ( .A1(n18366), .A2(n25891), .B1(n18338), .B2(n25890), .ZN(
        n13518) );
  AOI221_X2 U6061 ( .B1(n18351), .B2(n25887), .C1(n18342), .C2(n25885), .A(
        n13519), .ZN(n13508) );
  AOI221_X2 U6063 ( .B1(n18368), .B2(n25877), .C1(n18359), .C2(n25875), .A(
        n13522), .ZN(n13507) );
  OAI22_X2 U6064 ( .A1(n25873), .A2(n26673), .B1(n25871), .B2(n26689), .ZN(
        n13522) );
  NAND4_X2 U6065 ( .A1(n13525), .A2(n13526), .A3(n13527), .A4(n13528), .ZN(
        n13505) );
  AOI221_X2 U6066 ( .B1(n18340), .B2(n25869), .C1(n25868), .C2(n25519), .A(
        n13530), .ZN(n13528) );
  AOI221_X2 U6069 ( .B1(n25859), .B2(n25687), .C1(n25858), .C2(n25200), .A(
        n13536), .ZN(n13527) );
  OAI22_X2 U6070 ( .A1(n18371), .A2(n25855), .B1(n18343), .B2(n25854), .ZN(
        n13536) );
  AOI221_X2 U6073 ( .B1(n18363), .B2(n25851), .C1(n18354), .C2(n25850), .A(
        n13537), .ZN(n13526) );
  AOI221_X2 U6075 ( .B1(n18364), .B2(n25841), .C1(n18355), .C2(n25839), .A(
        n13538), .ZN(n13525) );
  OAI22_X2 U6076 ( .A1(n25837), .A2(n27137), .B1(n25835), .B2(n27201), .ZN(
        n13538) );
  NAND4_X2 U6079 ( .A1(n13544), .A2(n13545), .A3(n13546), .A4(n13547), .ZN(
        n13543) );
  AOI221_X2 U6080 ( .B1(n25905), .B2(n25030), .C1(n25903), .C2(n25518), .A(
        n13550), .ZN(n13547) );
  AOI221_X2 U6084 ( .B1(n25895), .B2(n25029), .C1(n25893), .C2(n25517), .A(
        n13555), .ZN(n13546) );
  OAI22_X2 U6085 ( .A1(n18329), .A2(n25891), .B1(n18301), .B2(n25889), .ZN(
        n13555) );
  AOI221_X2 U6088 ( .B1(n18314), .B2(n25888), .C1(n18305), .C2(n25886), .A(
        n13556), .ZN(n13545) );
  AOI221_X2 U6090 ( .B1(n18331), .B2(n25877), .C1(n18322), .C2(n25875), .A(
        n13559), .ZN(n13544) );
  OAI22_X2 U6091 ( .A1(n25873), .A2(n26674), .B1(n25872), .B2(n26690), .ZN(
        n13559) );
  NAND4_X2 U6092 ( .A1(n13562), .A2(n13563), .A3(n13564), .A4(n13565), .ZN(
        n13542) );
  AOI221_X2 U6093 ( .B1(n18303), .B2(n25870), .C1(n25867), .C2(n25516), .A(
        n13567), .ZN(n13565) );
  AOI221_X2 U6096 ( .B1(n25859), .B2(n25686), .C1(n25857), .C2(n25199), .A(
        n13573), .ZN(n13564) );
  OAI22_X2 U6097 ( .A1(n18334), .A2(n25855), .B1(n18306), .B2(n25853), .ZN(
        n13573) );
  AOI221_X2 U6100 ( .B1(n18326), .B2(n25851), .C1(n18317), .C2(n25849), .A(
        n13574), .ZN(n13563) );
  AOI221_X2 U6102 ( .B1(n18327), .B2(n25841), .C1(n18318), .C2(n25839), .A(
        n13575), .ZN(n13562) );
  OAI22_X2 U6103 ( .A1(n25837), .A2(n27138), .B1(n25835), .B2(n27202), .ZN(
        n13575) );
  OAI22_X2 U6104 ( .A1(n18298), .A2(n25907), .B1(n13578), .B2(n12153), .ZN(
        n23464) );
  NOR2_X2 U6105 ( .A1(n13579), .A2(n13580), .ZN(n13578) );
  NAND4_X2 U6106 ( .A1(n13581), .A2(n13582), .A3(n13583), .A4(n13584), .ZN(
        n13580) );
  AOI221_X2 U6107 ( .B1(n25905), .B2(n25685), .C1(n25904), .C2(n25198), .A(
        n13587), .ZN(n13584) );
  AOI221_X2 U6111 ( .B1(n25895), .B2(n25684), .C1(n25894), .C2(n25197), .A(
        n13592), .ZN(n13583) );
  OAI22_X2 U6112 ( .A1(n18292), .A2(n25892), .B1(n18264), .B2(n25890), .ZN(
        n13592) );
  AOI221_X2 U6115 ( .B1(n18277), .B2(n25887), .C1(n18268), .C2(n25885), .A(
        n13593), .ZN(n13582) );
  AOI221_X2 U6117 ( .B1(n18294), .B2(n25877), .C1(n18285), .C2(n25876), .A(
        n13596), .ZN(n13581) );
  OAI22_X2 U6118 ( .A1(n25873), .A2(n26675), .B1(n25871), .B2(n26691), .ZN(
        n13596) );
  NAND4_X2 U6119 ( .A1(n13599), .A2(n13600), .A3(n13601), .A4(n13602), .ZN(
        n13579) );
  AOI221_X2 U6120 ( .B1(n18266), .B2(n25870), .C1(n25867), .C2(n25515), .A(
        n13604), .ZN(n13602) );
  AOI221_X2 U6123 ( .B1(n25859), .B2(n25683), .C1(n25858), .C2(n25196), .A(
        n13610), .ZN(n13601) );
  OAI22_X2 U6124 ( .A1(n18297), .A2(n25856), .B1(n18269), .B2(n25854), .ZN(
        n13610) );
  AOI221_X2 U6127 ( .B1(n18289), .B2(n25851), .C1(n18280), .C2(n25850), .A(
        n13611), .ZN(n13600) );
  AOI221_X2 U6129 ( .B1(n18290), .B2(n25841), .C1(n18281), .C2(n25840), .A(
        n13612), .ZN(n13599) );
  OAI22_X2 U6130 ( .A1(n25837), .A2(n27139), .B1(n25835), .B2(n27203), .ZN(
        n13612) );
  OAI22_X2 U6131 ( .A1(n18261), .A2(n25909), .B1(n13615), .B2(n12153), .ZN(
        n23465) );
  NOR2_X2 U6132 ( .A1(n13616), .A2(n13617), .ZN(n13615) );
  NAND4_X2 U6133 ( .A1(n13618), .A2(n13619), .A3(n13620), .A4(n13621), .ZN(
        n13617) );
  AOI221_X2 U6134 ( .B1(n25906), .B2(n25682), .C1(n25904), .C2(n25195), .A(
        n13624), .ZN(n13621) );
  AOI221_X2 U6138 ( .B1(n25895), .B2(n25681), .C1(n25894), .C2(n25194), .A(
        n13629), .ZN(n13620) );
  OAI22_X2 U6139 ( .A1(n18255), .A2(n25892), .B1(n18227), .B2(n25890), .ZN(
        n13629) );
  AOI221_X2 U6142 ( .B1(n18240), .B2(n25887), .C1(n18231), .C2(n25885), .A(
        n13630), .ZN(n13619) );
  AOI221_X2 U6144 ( .B1(n18257), .B2(n25878), .C1(n18248), .C2(n25876), .A(
        n13633), .ZN(n13618) );
  OAI22_X2 U6145 ( .A1(n25873), .A2(n26676), .B1(n25871), .B2(n26692), .ZN(
        n13633) );
  NAND4_X2 U6146 ( .A1(n13636), .A2(n13637), .A3(n13638), .A4(n13639), .ZN(
        n13616) );
  AOI221_X2 U6147 ( .B1(n18229), .B2(n25869), .C1(n25868), .C2(n25514), .A(
        n13641), .ZN(n13639) );
  AOI221_X2 U6150 ( .B1(n25860), .B2(n25680), .C1(n25858), .C2(n25193), .A(
        n13647), .ZN(n13638) );
  OAI22_X2 U6151 ( .A1(n18260), .A2(n25856), .B1(n18232), .B2(n25853), .ZN(
        n13647) );
  AOI221_X2 U6154 ( .B1(n18252), .B2(n25852), .C1(n18243), .C2(n25850), .A(
        n13648), .ZN(n13637) );
  AOI221_X2 U6156 ( .B1(n18253), .B2(n25842), .C1(n18244), .C2(n25840), .A(
        n13649), .ZN(n13636) );
  OAI22_X2 U6157 ( .A1(n25837), .A2(n27140), .B1(n25835), .B2(n27204), .ZN(
        n13649) );
  OAI22_X2 U6158 ( .A1(n18224), .A2(n25907), .B1(n13652), .B2(n12153), .ZN(
        n23466) );
  NOR2_X2 U6159 ( .A1(n13653), .A2(n13654), .ZN(n13652) );
  NAND4_X2 U6160 ( .A1(n13655), .A2(n13656), .A3(n13657), .A4(n13658), .ZN(
        n13654) );
  AOI221_X2 U6161 ( .B1(n25906), .B2(n25679), .C1(n25903), .C2(n25192), .A(
        n13661), .ZN(n13658) );
  AOI221_X2 U6165 ( .B1(n25896), .B2(n25678), .C1(n25893), .C2(n25191), .A(
        n13666), .ZN(n13657) );
  OAI22_X2 U6166 ( .A1(n18218), .A2(n25892), .B1(n18190), .B2(n25890), .ZN(
        n13666) );
  AOI221_X2 U6169 ( .B1(n18203), .B2(n25887), .C1(n18194), .C2(n25885), .A(
        n13667), .ZN(n13656) );
  AOI221_X2 U6171 ( .B1(n18220), .B2(n25877), .C1(n18211), .C2(n25875), .A(
        n13670), .ZN(n13655) );
  OAI22_X2 U6172 ( .A1(n25873), .A2(n26677), .B1(n25871), .B2(n26693), .ZN(
        n13670) );
  NAND4_X2 U6173 ( .A1(n13673), .A2(n13674), .A3(n13675), .A4(n13676), .ZN(
        n13653) );
  AOI221_X2 U6174 ( .B1(n18192), .B2(n25869), .C1(n25868), .C2(n25513), .A(
        n13678), .ZN(n13676) );
  AOI221_X2 U6177 ( .B1(n25860), .B2(n25677), .C1(n25857), .C2(n25190), .A(
        n13684), .ZN(n13675) );
  OAI22_X2 U6178 ( .A1(n18223), .A2(n25856), .B1(n18195), .B2(n25853), .ZN(
        n13684) );
  AOI221_X2 U6181 ( .B1(n18215), .B2(n25851), .C1(n18206), .C2(n25849), .A(
        n13685), .ZN(n13674) );
  AOI221_X2 U6183 ( .B1(n18216), .B2(n25841), .C1(n18207), .C2(n25839), .A(
        n13686), .ZN(n13673) );
  OAI22_X2 U6184 ( .A1(n25838), .A2(n27141), .B1(n25835), .B2(n27205), .ZN(
        n13686) );
  OAI22_X2 U6185 ( .A1(n18187), .A2(n25909), .B1(n13689), .B2(n12153), .ZN(
        n23467) );
  NOR2_X2 U6186 ( .A1(n13690), .A2(n13691), .ZN(n13689) );
  NAND4_X2 U6187 ( .A1(n13692), .A2(n13693), .A3(n13694), .A4(n13695), .ZN(
        n13691) );
  AOI221_X2 U6188 ( .B1(n25906), .B2(n25676), .C1(n25903), .C2(n25189), .A(
        n13698), .ZN(n13695) );
  AOI221_X2 U6192 ( .B1(n25896), .B2(n25675), .C1(n25893), .C2(n25188), .A(
        n13703), .ZN(n13694) );
  OAI22_X2 U6193 ( .A1(n18181), .A2(n25892), .B1(n18153), .B2(n25890), .ZN(
        n13703) );
  AOI221_X2 U6196 ( .B1(n18166), .B2(n25887), .C1(n18157), .C2(n25885), .A(
        n13704), .ZN(n13693) );
  AOI221_X2 U6198 ( .B1(n18183), .B2(n25877), .C1(n18174), .C2(n25875), .A(
        n13707), .ZN(n13692) );
  OAI22_X2 U6199 ( .A1(n25873), .A2(n26678), .B1(n25871), .B2(n26694), .ZN(
        n13707) );
  NAND4_X2 U6200 ( .A1(n13710), .A2(n13711), .A3(n13712), .A4(n13713), .ZN(
        n13690) );
  AOI221_X2 U6201 ( .B1(n18155), .B2(n25869), .C1(n25867), .C2(n25512), .A(
        n13715), .ZN(n13713) );
  AOI221_X2 U6204 ( .B1(n25860), .B2(n25674), .C1(n25857), .C2(n25187), .A(
        n13721), .ZN(n13712) );
  OAI22_X2 U6205 ( .A1(n18186), .A2(n25856), .B1(n18158), .B2(n25854), .ZN(
        n13721) );
  AOI221_X2 U6208 ( .B1(n18178), .B2(n25851), .C1(n18169), .C2(n25850), .A(
        n13722), .ZN(n13711) );
  AOI221_X2 U6210 ( .B1(n18179), .B2(n25841), .C1(n18170), .C2(n25839), .A(
        n13723), .ZN(n13710) );
  OAI22_X2 U6211 ( .A1(n25838), .A2(n27142), .B1(n25835), .B2(n27206), .ZN(
        n13723) );
  NAND4_X2 U6214 ( .A1(n13729), .A2(n13730), .A3(n13731), .A4(n13732), .ZN(
        n13728) );
  AOI221_X2 U6215 ( .B1(n25906), .B2(n25028), .C1(n25903), .C2(n25511), .A(
        n13735), .ZN(n13732) );
  AOI221_X2 U6219 ( .B1(n25895), .B2(n25027), .C1(n25894), .C2(n25510), .A(
        n13740), .ZN(n13731) );
  OAI22_X2 U6220 ( .A1(n18144), .A2(n25892), .B1(n18116), .B2(n25889), .ZN(
        n13740) );
  AOI221_X2 U6223 ( .B1(n18129), .B2(n25887), .C1(n18120), .C2(n25885), .A(
        n13741), .ZN(n13730) );
  AOI221_X2 U6225 ( .B1(n18146), .B2(n25878), .C1(n18137), .C2(n25875), .A(
        n13744), .ZN(n13729) );
  OAI22_X2 U6226 ( .A1(n25874), .A2(n26727), .B1(n25871), .B2(n26743), .ZN(
        n13744) );
  NAND4_X2 U6227 ( .A1(n13747), .A2(n13748), .A3(n13749), .A4(n13750), .ZN(
        n13727) );
  AOI221_X2 U6228 ( .B1(n18118), .B2(n25869), .C1(n25867), .C2(n25509), .A(
        n13752), .ZN(n13750) );
  AOI221_X2 U6231 ( .B1(n25860), .B2(n25673), .C1(n25857), .C2(n25186), .A(
        n13758), .ZN(n13749) );
  OAI22_X2 U6232 ( .A1(n18149), .A2(n25856), .B1(n18121), .B2(n25854), .ZN(
        n13758) );
  AOI221_X2 U6235 ( .B1(n18141), .B2(n25852), .C1(n18132), .C2(n25849), .A(
        n13759), .ZN(n13748) );
  AOI221_X2 U6237 ( .B1(n18142), .B2(n25842), .C1(n18133), .C2(n25839), .A(
        n13760), .ZN(n13747) );
  OAI22_X2 U6238 ( .A1(n25837), .A2(n27111), .B1(n25835), .B2(n27175), .ZN(
        n13760) );
  NAND4_X2 U6241 ( .A1(n13766), .A2(n13767), .A3(n13768), .A4(n13769), .ZN(
        n13765) );
  AOI221_X2 U6242 ( .B1(n25906), .B2(n25026), .C1(n25904), .C2(n25508), .A(
        n13772), .ZN(n13769) );
  AOI221_X2 U6246 ( .B1(n25896), .B2(n25025), .C1(n25894), .C2(n25507), .A(
        n13777), .ZN(n13768) );
  OAI22_X2 U6247 ( .A1(n18107), .A2(n25892), .B1(n18079), .B2(n25889), .ZN(
        n13777) );
  AOI221_X2 U6250 ( .B1(n18092), .B2(n25887), .C1(n18083), .C2(n25885), .A(
        n13778), .ZN(n13767) );
  AOI221_X2 U6252 ( .B1(n18109), .B2(n25877), .C1(n18100), .C2(n25876), .A(
        n13781), .ZN(n13766) );
  OAI22_X2 U6253 ( .A1(n25873), .A2(n26728), .B1(n25871), .B2(n26744), .ZN(
        n13781) );
  NAND4_X2 U6254 ( .A1(n13784), .A2(n13785), .A3(n13786), .A4(n13787), .ZN(
        n13764) );
  AOI221_X2 U6255 ( .B1(n18081), .B2(n25869), .C1(n25868), .C2(n25506), .A(
        n13789), .ZN(n13787) );
  AOI221_X2 U6258 ( .B1(n25860), .B2(n25672), .C1(n25858), .C2(n25185), .A(
        n13795), .ZN(n13786) );
  OAI22_X2 U6259 ( .A1(n18112), .A2(n25856), .B1(n18084), .B2(n25853), .ZN(
        n13795) );
  AOI221_X2 U6262 ( .B1(n18104), .B2(n25851), .C1(n18095), .C2(n25850), .A(
        n13796), .ZN(n13785) );
  AOI221_X2 U6264 ( .B1(n18105), .B2(n25841), .C1(n18096), .C2(n25840), .A(
        n13797), .ZN(n13784) );
  OAI22_X2 U6265 ( .A1(n25838), .A2(n27112), .B1(n25835), .B2(n27176), .ZN(
        n13797) );
  NAND4_X2 U6268 ( .A1(n13803), .A2(n13804), .A3(n13805), .A4(n13806), .ZN(
        n13802) );
  AOI221_X2 U6269 ( .B1(n25906), .B2(n25024), .C1(n25904), .C2(n25505), .A(
        n13809), .ZN(n13806) );
  AOI221_X2 U6273 ( .B1(n25895), .B2(n25023), .C1(n25893), .C2(n25504), .A(
        n13814), .ZN(n13805) );
  OAI22_X2 U6274 ( .A1(n18070), .A2(n25892), .B1(n18042), .B2(n25890), .ZN(
        n13814) );
  AOI221_X2 U6277 ( .B1(n18055), .B2(n25887), .C1(n18046), .C2(n25885), .A(
        n13815), .ZN(n13804) );
  AOI221_X2 U6279 ( .B1(n18072), .B2(n25878), .C1(n18063), .C2(n25875), .A(
        n13818), .ZN(n13803) );
  OAI22_X2 U6280 ( .A1(n25874), .A2(n26729), .B1(n25871), .B2(n26745), .ZN(
        n13818) );
  NAND4_X2 U6281 ( .A1(n13821), .A2(n13822), .A3(n13823), .A4(n13824), .ZN(
        n13801) );
  AOI221_X2 U6282 ( .B1(n18044), .B2(n25869), .C1(n25867), .C2(n25503), .A(
        n13826), .ZN(n13824) );
  AOI221_X2 U6285 ( .B1(n25860), .B2(n25671), .C1(n25858), .C2(n25184), .A(
        n13832), .ZN(n13823) );
  OAI22_X2 U6286 ( .A1(n18075), .A2(n25856), .B1(n18047), .B2(n25854), .ZN(
        n13832) );
  AOI221_X2 U6289 ( .B1(n18067), .B2(n25852), .C1(n18058), .C2(n25850), .A(
        n13833), .ZN(n13822) );
  AOI221_X2 U6291 ( .B1(n18068), .B2(n25842), .C1(n18059), .C2(n25839), .A(
        n13834), .ZN(n13821) );
  OAI22_X2 U6292 ( .A1(n25837), .A2(n27113), .B1(n25835), .B2(n27177), .ZN(
        n13834) );
  NAND4_X2 U6295 ( .A1(n13840), .A2(n13841), .A3(n13842), .A4(n13843), .ZN(
        n13839) );
  AOI221_X2 U6296 ( .B1(n25906), .B2(n25022), .C1(n25903), .C2(n25502), .A(
        n13846), .ZN(n13843) );
  AOI221_X2 U6300 ( .B1(n25895), .B2(n25021), .C1(n25894), .C2(n25501), .A(
        n13851), .ZN(n13842) );
  OAI22_X2 U6301 ( .A1(n18033), .A2(n25892), .B1(n18005), .B2(n25889), .ZN(
        n13851) );
  AOI221_X2 U6304 ( .B1(n18018), .B2(n25887), .C1(n18009), .C2(n25885), .A(
        n13852), .ZN(n13841) );
  AOI221_X2 U6306 ( .B1(n18035), .B2(n25877), .C1(n18026), .C2(n25875), .A(
        n13855), .ZN(n13840) );
  OAI22_X2 U6307 ( .A1(n25873), .A2(n26730), .B1(n25871), .B2(n26746), .ZN(
        n13855) );
  NAND4_X2 U6308 ( .A1(n13858), .A2(n13859), .A3(n13860), .A4(n13861), .ZN(
        n13838) );
  AOI221_X2 U6309 ( .B1(n18007), .B2(n25869), .C1(n25867), .C2(n25500), .A(
        n13863), .ZN(n13861) );
  AOI221_X2 U6312 ( .B1(n25860), .B2(n25670), .C1(n25857), .C2(n25183), .A(
        n13869), .ZN(n13860) );
  OAI22_X2 U6313 ( .A1(n18038), .A2(n25856), .B1(n18010), .B2(n25853), .ZN(
        n13869) );
  AOI221_X2 U6316 ( .B1(n18030), .B2(n25851), .C1(n18021), .C2(n25849), .A(
        n13870), .ZN(n13859) );
  AOI221_X2 U6318 ( .B1(n18031), .B2(n25841), .C1(n18022), .C2(n25839), .A(
        n13871), .ZN(n13858) );
  OAI22_X2 U6319 ( .A1(n25838), .A2(n27114), .B1(n25835), .B2(n27178), .ZN(
        n13871) );
  NAND4_X2 U6322 ( .A1(n13877), .A2(n13878), .A3(n13879), .A4(n13880), .ZN(
        n13876) );
  AOI221_X2 U6323 ( .B1(n25906), .B2(n25020), .C1(n25904), .C2(n25499), .A(
        n13883), .ZN(n13880) );
  AOI221_X2 U6327 ( .B1(n25896), .B2(n25019), .C1(n25893), .C2(n25498), .A(
        n13888), .ZN(n13879) );
  OAI22_X2 U6328 ( .A1(n17996), .A2(n25892), .B1(n17968), .B2(n25889), .ZN(
        n13888) );
  AOI221_X2 U6331 ( .B1(n17981), .B2(n25887), .C1(n17972), .C2(n25885), .A(
        n13889), .ZN(n13878) );
  AOI221_X2 U6333 ( .B1(n17998), .B2(n25878), .C1(n17989), .C2(n25876), .A(
        n13892), .ZN(n13877) );
  OAI22_X2 U6334 ( .A1(n25874), .A2(n26731), .B1(n25871), .B2(n26747), .ZN(
        n13892) );
  NAND4_X2 U6335 ( .A1(n13895), .A2(n13896), .A3(n13897), .A4(n13898), .ZN(
        n13875) );
  AOI221_X2 U6336 ( .B1(n17970), .B2(n25869), .C1(n25868), .C2(n25497), .A(
        n13900), .ZN(n13898) );
  AOI221_X2 U6339 ( .B1(n25860), .B2(n25669), .C1(n25858), .C2(n25182), .A(
        n13906), .ZN(n13897) );
  OAI22_X2 U6340 ( .A1(n18001), .A2(n25856), .B1(n17973), .B2(n25853), .ZN(
        n13906) );
  AOI221_X2 U6343 ( .B1(n17993), .B2(n25852), .C1(n17984), .C2(n25850), .A(
        n13907), .ZN(n13896) );
  AOI221_X2 U6345 ( .B1(n17994), .B2(n25842), .C1(n17985), .C2(n25840), .A(
        n13908), .ZN(n13895) );
  OAI22_X2 U6346 ( .A1(n25837), .A2(n27115), .B1(n25835), .B2(n27179), .ZN(
        n13908) );
  NAND4_X2 U6349 ( .A1(n13914), .A2(n13915), .A3(n13916), .A4(n13917), .ZN(
        n13913) );
  AOI221_X2 U6350 ( .B1(n25906), .B2(n25018), .C1(n25903), .C2(n25496), .A(
        n13920), .ZN(n13917) );
  AOI221_X2 U6354 ( .B1(n25896), .B2(n25017), .C1(n25893), .C2(n25495), .A(
        n13925), .ZN(n13916) );
  OAI22_X2 U6355 ( .A1(n17959), .A2(n25892), .B1(n17931), .B2(n25889), .ZN(
        n13925) );
  AOI221_X2 U6358 ( .B1(n17944), .B2(n25887), .C1(n17935), .C2(n25885), .A(
        n13926), .ZN(n13915) );
  AOI221_X2 U6360 ( .B1(n17961), .B2(n25877), .C1(n17952), .C2(n25876), .A(
        n13929), .ZN(n13914) );
  OAI22_X2 U6361 ( .A1(n25873), .A2(n26732), .B1(n25871), .B2(n26748), .ZN(
        n13929) );
  NAND4_X2 U6362 ( .A1(n13932), .A2(n13933), .A3(n13934), .A4(n13935), .ZN(
        n13912) );
  AOI221_X2 U6363 ( .B1(n17933), .B2(n25869), .C1(n25868), .C2(n25494), .A(
        n13937), .ZN(n13935) );
  AOI221_X2 U6366 ( .B1(n25860), .B2(n25668), .C1(n25857), .C2(n25181), .A(
        n13943), .ZN(n13934) );
  OAI22_X2 U6367 ( .A1(n17964), .A2(n25856), .B1(n17936), .B2(n25853), .ZN(
        n13943) );
  AOI221_X2 U6370 ( .B1(n17956), .B2(n25851), .C1(n17947), .C2(n25849), .A(
        n13944), .ZN(n13933) );
  AOI221_X2 U6372 ( .B1(n17957), .B2(n25841), .C1(n17948), .C2(n25840), .A(
        n13945), .ZN(n13932) );
  OAI22_X2 U6373 ( .A1(n25838), .A2(n27116), .B1(n25835), .B2(n27180), .ZN(
        n13945) );
  NAND4_X2 U6376 ( .A1(n13951), .A2(n13952), .A3(n13953), .A4(n13954), .ZN(
        n13950) );
  AOI221_X2 U6377 ( .B1(n25906), .B2(n25016), .C1(n25903), .C2(n25493), .A(
        n13957), .ZN(n13954) );
  AOI221_X2 U6381 ( .B1(n25895), .B2(n25015), .C1(n25894), .C2(n25492), .A(
        n13962), .ZN(n13953) );
  OAI22_X2 U6382 ( .A1(n17922), .A2(n25892), .B1(n17894), .B2(n25890), .ZN(
        n13962) );
  AOI221_X2 U6385 ( .B1(n17907), .B2(n25887), .C1(n17898), .C2(n25885), .A(
        n13963), .ZN(n13952) );
  AOI221_X2 U6387 ( .B1(n17924), .B2(n25878), .C1(n17915), .C2(n25875), .A(
        n13966), .ZN(n13951) );
  OAI22_X2 U6388 ( .A1(n25874), .A2(n26733), .B1(n25871), .B2(n26749), .ZN(
        n13966) );
  NAND4_X2 U6389 ( .A1(n13969), .A2(n13970), .A3(n13971), .A4(n13972), .ZN(
        n13949) );
  AOI221_X2 U6390 ( .B1(n17896), .B2(n25869), .C1(n25867), .C2(n25491), .A(
        n13974), .ZN(n13972) );
  AOI221_X2 U6393 ( .B1(n25860), .B2(n25667), .C1(n25857), .C2(n25180), .A(
        n13980), .ZN(n13971) );
  OAI22_X2 U6394 ( .A1(n17927), .A2(n25856), .B1(n17899), .B2(n25853), .ZN(
        n13980) );
  AOI221_X2 U6397 ( .B1(n17919), .B2(n25852), .C1(n17910), .C2(n25849), .A(
        n13981), .ZN(n13970) );
  AOI221_X2 U6399 ( .B1(n17920), .B2(n25842), .C1(n17911), .C2(n25839), .A(
        n13982), .ZN(n13969) );
  OAI22_X2 U6400 ( .A1(n25837), .A2(n27117), .B1(n25835), .B2(n27181), .ZN(
        n13982) );
  NAND4_X2 U6403 ( .A1(n13988), .A2(n13989), .A3(n13990), .A4(n13991), .ZN(
        n13987) );
  AOI221_X2 U6404 ( .B1(n25906), .B2(n25014), .C1(n25904), .C2(n25490), .A(
        n13994), .ZN(n13991) );
  AOI221_X2 U6408 ( .B1(n25896), .B2(n25013), .C1(n25894), .C2(n25489), .A(
        n13999), .ZN(n13990) );
  OAI22_X2 U6409 ( .A1(n17885), .A2(n25892), .B1(n17857), .B2(n25889), .ZN(
        n13999) );
  AOI221_X2 U6412 ( .B1(n17870), .B2(n25887), .C1(n17861), .C2(n25885), .A(
        n14000), .ZN(n13989) );
  AOI221_X2 U6414 ( .B1(n17887), .B2(n25877), .C1(n17878), .C2(n25876), .A(
        n14003), .ZN(n13988) );
  OAI22_X2 U6415 ( .A1(n25873), .A2(n26734), .B1(n25871), .B2(n26750), .ZN(
        n14003) );
  NAND4_X2 U6416 ( .A1(n14006), .A2(n14007), .A3(n14008), .A4(n14009), .ZN(
        n13986) );
  AOI221_X2 U6417 ( .B1(n17859), .B2(n25869), .C1(n25868), .C2(n25488), .A(
        n14011), .ZN(n14009) );
  AOI221_X2 U6420 ( .B1(n25860), .B2(n25666), .C1(n25858), .C2(n25179), .A(
        n14017), .ZN(n14008) );
  OAI22_X2 U6421 ( .A1(n17890), .A2(n25856), .B1(n17862), .B2(n25853), .ZN(
        n14017) );
  AOI221_X2 U6424 ( .B1(n17882), .B2(n25851), .C1(n17873), .C2(n25850), .A(
        n14018), .ZN(n14007) );
  AOI221_X2 U6426 ( .B1(n17883), .B2(n25841), .C1(n17874), .C2(n25840), .A(
        n14019), .ZN(n14006) );
  OAI22_X2 U6427 ( .A1(n25838), .A2(n27118), .B1(n25835), .B2(n27182), .ZN(
        n14019) );
  NAND4_X2 U6430 ( .A1(n14025), .A2(n14026), .A3(n14027), .A4(n14028), .ZN(
        n14024) );
  AOI221_X2 U6431 ( .B1(n25906), .B2(n25012), .C1(n25904), .C2(n25487), .A(
        n14031), .ZN(n14028) );
  AOI221_X2 U6435 ( .B1(n25896), .B2(n25011), .C1(n25893), .C2(n25486), .A(
        n14036), .ZN(n14027) );
  OAI22_X2 U6436 ( .A1(n17848), .A2(n25891), .B1(n17820), .B2(n25889), .ZN(
        n14036) );
  AOI221_X2 U6439 ( .B1(n17833), .B2(n25887), .C1(n17824), .C2(n25885), .A(
        n14037), .ZN(n14026) );
  AOI221_X2 U6441 ( .B1(n17850), .B2(n25878), .C1(n17841), .C2(n25876), .A(
        n14040), .ZN(n14025) );
  OAI22_X2 U6442 ( .A1(n25874), .A2(n26735), .B1(n25871), .B2(n26751), .ZN(
        n14040) );
  NAND4_X2 U6443 ( .A1(n14043), .A2(n14044), .A3(n14045), .A4(n14046), .ZN(
        n14023) );
  AOI221_X2 U6444 ( .B1(n17822), .B2(n25869), .C1(n25867), .C2(n25485), .A(
        n14048), .ZN(n14046) );
  AOI221_X2 U6447 ( .B1(n25860), .B2(n25665), .C1(n25858), .C2(n25178), .A(
        n14054), .ZN(n14045) );
  OAI22_X2 U6448 ( .A1(n17853), .A2(n25856), .B1(n17825), .B2(n25853), .ZN(
        n14054) );
  AOI221_X2 U6451 ( .B1(n17845), .B2(n25852), .C1(n17836), .C2(n25850), .A(
        n14055), .ZN(n14044) );
  AOI221_X2 U6453 ( .B1(n17846), .B2(n25842), .C1(n17837), .C2(n25840), .A(
        n14056), .ZN(n14043) );
  OAI22_X2 U6454 ( .A1(n25838), .A2(n27119), .B1(n25835), .B2(n27183), .ZN(
        n14056) );
  NAND4_X2 U6457 ( .A1(n14062), .A2(n14063), .A3(n14064), .A4(n14065), .ZN(
        n14061) );
  AOI221_X2 U6458 ( .B1(n25906), .B2(n25010), .C1(n25903), .C2(n25484), .A(
        n14068), .ZN(n14065) );
  AOI221_X2 U6462 ( .B1(n25895), .B2(n25009), .C1(n25894), .C2(n25483), .A(
        n14073), .ZN(n14064) );
  OAI22_X2 U6463 ( .A1(n17811), .A2(n25892), .B1(n17783), .B2(n25889), .ZN(
        n14073) );
  AOI221_X2 U6466 ( .B1(n17796), .B2(n25887), .C1(n17787), .C2(n25885), .A(
        n14074), .ZN(n14063) );
  AOI221_X2 U6468 ( .B1(n17813), .B2(n25877), .C1(n17804), .C2(n25875), .A(
        n14077), .ZN(n14062) );
  OAI22_X2 U6469 ( .A1(n25873), .A2(n26736), .B1(n25871), .B2(n26752), .ZN(
        n14077) );
  NAND4_X2 U6470 ( .A1(n14080), .A2(n14081), .A3(n14082), .A4(n14083), .ZN(
        n14060) );
  AOI221_X2 U6471 ( .B1(n17785), .B2(n25869), .C1(n25867), .C2(n25482), .A(
        n14085), .ZN(n14083) );
  AOI221_X2 U6474 ( .B1(n25860), .B2(n25664), .C1(n25857), .C2(n25177), .A(
        n14091), .ZN(n14082) );
  OAI22_X2 U6475 ( .A1(n17816), .A2(n25855), .B1(n17788), .B2(n25853), .ZN(
        n14091) );
  AOI221_X2 U6478 ( .B1(n17808), .B2(n25851), .C1(n17799), .C2(n25849), .A(
        n14092), .ZN(n14081) );
  AOI221_X2 U6480 ( .B1(n17809), .B2(n25841), .C1(n17800), .C2(n25839), .A(
        n14093), .ZN(n14080) );
  OAI22_X2 U6481 ( .A1(n25838), .A2(n27120), .B1(n25836), .B2(n27184), .ZN(
        n14093) );
  NAND4_X2 U6484 ( .A1(n14099), .A2(n14100), .A3(n14101), .A4(n14102), .ZN(
        n14098) );
  AOI221_X2 U6485 ( .B1(n25905), .B2(n25008), .C1(n25903), .C2(n25481), .A(
        n14105), .ZN(n14102) );
  AOI221_X2 U6489 ( .B1(n25896), .B2(n25007), .C1(n25893), .C2(n25480), .A(
        n14110), .ZN(n14101) );
  OAI22_X2 U6490 ( .A1(n17774), .A2(n25891), .B1(n17746), .B2(n25889), .ZN(
        n14110) );
  AOI221_X2 U6493 ( .B1(n17759), .B2(n25888), .C1(n17750), .C2(n25886), .A(
        n14111), .ZN(n14100) );
  AOI221_X2 U6495 ( .B1(n17776), .B2(n25878), .C1(n17767), .C2(n25875), .A(
        n14114), .ZN(n14099) );
  OAI22_X2 U6496 ( .A1(n25874), .A2(n26737), .B1(n25872), .B2(n26753), .ZN(
        n14114) );
  NAND4_X2 U6497 ( .A1(n14117), .A2(n14118), .A3(n14119), .A4(n14120), .ZN(
        n14097) );
  AOI221_X2 U6498 ( .B1(n17748), .B2(n25870), .C1(n25867), .C2(n25479), .A(
        n14122), .ZN(n14120) );
  AOI221_X2 U6501 ( .B1(n25859), .B2(n25663), .C1(n25857), .C2(n25176), .A(
        n14128), .ZN(n14119) );
  OAI22_X2 U6502 ( .A1(n17779), .A2(n25856), .B1(n17751), .B2(n25853), .ZN(
        n14128) );
  AOI221_X2 U6505 ( .B1(n17771), .B2(n25852), .C1(n17762), .C2(n25849), .A(
        n14129), .ZN(n14118) );
  AOI221_X2 U6507 ( .B1(n17772), .B2(n25842), .C1(n17763), .C2(n25839), .A(
        n14130), .ZN(n14117) );
  OAI22_X2 U6508 ( .A1(n25838), .A2(n27121), .B1(n25835), .B2(n27185), .ZN(
        n14130) );
  NAND4_X2 U6511 ( .A1(n14136), .A2(n14137), .A3(n14138), .A4(n14139), .ZN(
        n14135) );
  AOI221_X2 U6512 ( .B1(n25906), .B2(n25006), .C1(n25903), .C2(n25478), .A(
        n14142), .ZN(n14139) );
  AOI221_X2 U6516 ( .B1(n25896), .B2(n25005), .C1(n25893), .C2(n25477), .A(
        n14147), .ZN(n14138) );
  OAI22_X2 U6517 ( .A1(n17737), .A2(n25892), .B1(n17709), .B2(n25889), .ZN(
        n14147) );
  AOI221_X2 U6520 ( .B1(n17722), .B2(n25888), .C1(n17713), .C2(n25886), .A(
        n14148), .ZN(n14137) );
  AOI221_X2 U6522 ( .B1(n17739), .B2(n25878), .C1(n17730), .C2(n25875), .A(
        n14151), .ZN(n14136) );
  OAI22_X2 U6523 ( .A1(n25873), .A2(n26738), .B1(n25871), .B2(n26754), .ZN(
        n14151) );
  NAND4_X2 U6524 ( .A1(n14154), .A2(n14155), .A3(n14156), .A4(n14157), .ZN(
        n14134) );
  AOI221_X2 U6525 ( .B1(n17711), .B2(n25870), .C1(n25867), .C2(n25476), .A(
        n14159), .ZN(n14157) );
  AOI221_X2 U6528 ( .B1(n25860), .B2(n25662), .C1(n25857), .C2(n25175), .A(
        n14165), .ZN(n14156) );
  OAI22_X2 U6529 ( .A1(n17742), .A2(n25855), .B1(n17714), .B2(n25853), .ZN(
        n14165) );
  AOI221_X2 U6532 ( .B1(n17734), .B2(n25852), .C1(n17725), .C2(n25849), .A(
        n14166), .ZN(n14155) );
  AOI221_X2 U6534 ( .B1(n17735), .B2(n25842), .C1(n17726), .C2(n25839), .A(
        n14167), .ZN(n14154) );
  OAI22_X2 U6535 ( .A1(n25838), .A2(n27122), .B1(n25836), .B2(n27186), .ZN(
        n14167) );
  OAI22_X2 U6536 ( .A1(n17706), .A2(n25907), .B1(n14170), .B2(n12153), .ZN(
        n23480) );
  NOR2_X2 U6537 ( .A1(n14171), .A2(n14172), .ZN(n14170) );
  NAND4_X2 U6538 ( .A1(n14173), .A2(n14174), .A3(n14175), .A4(n14176), .ZN(
        n14172) );
  AOI221_X2 U6539 ( .B1(n25905), .B2(n25661), .C1(n25903), .C2(n25174), .A(
        n14179), .ZN(n14176) );
  AOI221_X2 U6543 ( .B1(n25896), .B2(n25660), .C1(n25893), .C2(n25173), .A(
        n14184), .ZN(n14175) );
  OAI22_X2 U6544 ( .A1(n17700), .A2(n25891), .B1(n17672), .B2(n25889), .ZN(
        n14184) );
  AOI221_X2 U6547 ( .B1(n17685), .B2(n25888), .C1(n17676), .C2(n25886), .A(
        n14185), .ZN(n14174) );
  AOI221_X2 U6549 ( .B1(n17702), .B2(n25878), .C1(n17693), .C2(n25875), .A(
        n14188), .ZN(n14173) );
  OAI22_X2 U6550 ( .A1(n25873), .A2(n26739), .B1(n25871), .B2(n26755), .ZN(
        n14188) );
  NAND4_X2 U6551 ( .A1(n14191), .A2(n14192), .A3(n14193), .A4(n14194), .ZN(
        n14171) );
  AOI221_X2 U6552 ( .B1(n17674), .B2(n25870), .C1(n25867), .C2(n25475), .A(
        n14196), .ZN(n14194) );
  AOI221_X2 U6555 ( .B1(n25860), .B2(n25659), .C1(n25857), .C2(n25172), .A(
        n14202), .ZN(n14193) );
  OAI22_X2 U6556 ( .A1(n17705), .A2(n25855), .B1(n17677), .B2(n25853), .ZN(
        n14202) );
  AOI221_X2 U6559 ( .B1(n17697), .B2(n25852), .C1(n17688), .C2(n25849), .A(
        n14203), .ZN(n14192) );
  AOI221_X2 U6561 ( .B1(n17698), .B2(n25842), .C1(n17689), .C2(n25839), .A(
        n14204), .ZN(n14191) );
  OAI22_X2 U6562 ( .A1(n25838), .A2(n27123), .B1(n25835), .B2(n27187), .ZN(
        n14204) );
  OAI22_X2 U6563 ( .A1(n17669), .A2(n25909), .B1(n14207), .B2(n12153), .ZN(
        n23481) );
  NOR2_X2 U6564 ( .A1(n14208), .A2(n14209), .ZN(n14207) );
  NAND4_X2 U6565 ( .A1(n14210), .A2(n14211), .A3(n14212), .A4(n14213), .ZN(
        n14209) );
  AOI221_X2 U6566 ( .B1(n25906), .B2(n25658), .C1(n25903), .C2(n25171), .A(
        n14216), .ZN(n14213) );
  AOI221_X2 U6570 ( .B1(n25896), .B2(n25657), .C1(n25893), .C2(n25170), .A(
        n14221), .ZN(n14212) );
  OAI22_X2 U6571 ( .A1(n17663), .A2(n25891), .B1(n17635), .B2(n25889), .ZN(
        n14221) );
  AOI221_X2 U6574 ( .B1(n17648), .B2(n25888), .C1(n17639), .C2(n25886), .A(
        n14222), .ZN(n14211) );
  AOI221_X2 U6576 ( .B1(n17665), .B2(n25878), .C1(n17656), .C2(n25875), .A(
        n14225), .ZN(n14210) );
  OAI22_X2 U6577 ( .A1(n25874), .A2(n26740), .B1(n25871), .B2(n26756), .ZN(
        n14225) );
  NAND4_X2 U6578 ( .A1(n14228), .A2(n14229), .A3(n14230), .A4(n14231), .ZN(
        n14208) );
  AOI221_X2 U6579 ( .B1(n17637), .B2(n25870), .C1(n25867), .C2(n25474), .A(
        n14233), .ZN(n14231) );
  AOI221_X2 U6582 ( .B1(n25859), .B2(n25656), .C1(n25857), .C2(n25169), .A(
        n14239), .ZN(n14230) );
  OAI22_X2 U6583 ( .A1(n17668), .A2(n25855), .B1(n17640), .B2(n25853), .ZN(
        n14239) );
  AOI221_X2 U6586 ( .B1(n17660), .B2(n25852), .C1(n17651), .C2(n25849), .A(
        n14240), .ZN(n14229) );
  AOI221_X2 U6588 ( .B1(n17661), .B2(n25842), .C1(n17652), .C2(n25839), .A(
        n14241), .ZN(n14228) );
  OAI22_X2 U6589 ( .A1(n25838), .A2(n27124), .B1(n25836), .B2(n27188), .ZN(
        n14241) );
  OAI22_X2 U6590 ( .A1(n17632), .A2(n25907), .B1(n14244), .B2(n12153), .ZN(
        n23482) );
  NOR2_X2 U6591 ( .A1(n14245), .A2(n14246), .ZN(n14244) );
  NAND4_X2 U6592 ( .A1(n14247), .A2(n14248), .A3(n14249), .A4(n14250), .ZN(
        n14246) );
  AOI221_X2 U6593 ( .B1(n25906), .B2(n25655), .C1(n25903), .C2(n25168), .A(
        n14253), .ZN(n14250) );
  AOI221_X2 U6597 ( .B1(n25896), .B2(n25654), .C1(n25893), .C2(n25167), .A(
        n14258), .ZN(n14249) );
  OAI22_X2 U6598 ( .A1(n17626), .A2(n25892), .B1(n17598), .B2(n25889), .ZN(
        n14258) );
  AOI221_X2 U6601 ( .B1(n17611), .B2(n25888), .C1(n17602), .C2(n25886), .A(
        n14259), .ZN(n14248) );
  AOI221_X2 U6603 ( .B1(n17628), .B2(n25878), .C1(n17619), .C2(n25875), .A(
        n14262), .ZN(n14247) );
  OAI22_X2 U6604 ( .A1(n25874), .A2(n26741), .B1(n25872), .B2(n26757), .ZN(
        n14262) );
  NAND4_X2 U6605 ( .A1(n14265), .A2(n14266), .A3(n14267), .A4(n14268), .ZN(
        n14245) );
  AOI221_X2 U6606 ( .B1(n17600), .B2(n25870), .C1(n25867), .C2(n25473), .A(
        n14270), .ZN(n14268) );
  AOI221_X2 U6609 ( .B1(n25859), .B2(n25653), .C1(n25857), .C2(n25166), .A(
        n14276), .ZN(n14267) );
  OAI22_X2 U6610 ( .A1(n17631), .A2(n25856), .B1(n17603), .B2(n25853), .ZN(
        n14276) );
  AOI221_X2 U6613 ( .B1(n17623), .B2(n25852), .C1(n17614), .C2(n25849), .A(
        n14277), .ZN(n14266) );
  AOI221_X2 U6615 ( .B1(n17624), .B2(n25842), .C1(n17615), .C2(n25839), .A(
        n14278), .ZN(n14265) );
  OAI22_X2 U6616 ( .A1(n25838), .A2(n27125), .B1(n25836), .B2(n27189), .ZN(
        n14278) );
  OAI22_X2 U6617 ( .A1(n17595), .A2(n25909), .B1(n14281), .B2(n12153), .ZN(
        n23483) );
  NOR2_X2 U6618 ( .A1(n14282), .A2(n14283), .ZN(n14281) );
  NAND4_X2 U6619 ( .A1(n14284), .A2(n14285), .A3(n14286), .A4(n14287), .ZN(
        n14283) );
  AOI221_X2 U6620 ( .B1(n25905), .B2(n25652), .C1(n25903), .C2(n25165), .A(
        n14290), .ZN(n14287) );
  AOI221_X2 U6624 ( .B1(n25896), .B2(n25651), .C1(n25893), .C2(n25164), .A(
        n14295), .ZN(n14286) );
  OAI22_X2 U6625 ( .A1(n17589), .A2(n25892), .B1(n17561), .B2(n25889), .ZN(
        n14295) );
  AOI221_X2 U6628 ( .B1(n17574), .B2(n25888), .C1(n17565), .C2(n25886), .A(
        n14296), .ZN(n14285) );
  AOI221_X2 U6630 ( .B1(n17591), .B2(n25878), .C1(n17582), .C2(n25875), .A(
        n14299), .ZN(n14284) );
  OAI22_X2 U6631 ( .A1(n25874), .A2(n26742), .B1(n25872), .B2(n26758), .ZN(
        n14299) );
  NAND4_X2 U6632 ( .A1(n14302), .A2(n14303), .A3(n14304), .A4(n14305), .ZN(
        n14282) );
  AOI221_X2 U6633 ( .B1(n17563), .B2(n25870), .C1(n25867), .C2(n25472), .A(
        n14307), .ZN(n14305) );
  AOI221_X2 U6636 ( .B1(n25860), .B2(n25650), .C1(n25857), .C2(n25163), .A(
        n14313), .ZN(n14304) );
  OAI22_X2 U6637 ( .A1(n17594), .A2(n25856), .B1(n17566), .B2(n25853), .ZN(
        n14313) );
  AOI221_X2 U6640 ( .B1(n17586), .B2(n25852), .C1(n17577), .C2(n25849), .A(
        n14314), .ZN(n14303) );
  AOI221_X2 U6642 ( .B1(n17587), .B2(n25842), .C1(n17578), .C2(n25839), .A(
        n14315), .ZN(n14302) );
  OAI22_X2 U6643 ( .A1(n25838), .A2(n27126), .B1(n25835), .B2(n27190), .ZN(
        n14315) );
  NAND4_X2 U6646 ( .A1(n14321), .A2(n14322), .A3(n14323), .A4(n14324), .ZN(
        n14320) );
  AOI221_X2 U6647 ( .B1(n25905), .B2(n25004), .C1(n25903), .C2(n25471), .A(
        n14327), .ZN(n14324) );
  AOI221_X2 U6651 ( .B1(n25896), .B2(n25003), .C1(n25893), .C2(n25470), .A(
        n14332), .ZN(n14323) );
  OAI22_X2 U6652 ( .A1(n17552), .A2(n25892), .B1(n17524), .B2(n25889), .ZN(
        n14332) );
  AOI221_X2 U6655 ( .B1(n17537), .B2(n25888), .C1(n17528), .C2(n25886), .A(
        n14333), .ZN(n14322) );
  AOI221_X2 U6657 ( .B1(n17554), .B2(n25878), .C1(n17545), .C2(n25875), .A(
        n14336), .ZN(n14321) );
  OAI22_X2 U6658 ( .A1(n25873), .A2(n26519), .B1(n25872), .B2(n26615), .ZN(
        n14336) );
  NAND4_X2 U6659 ( .A1(n14339), .A2(n14340), .A3(n14341), .A4(n14342), .ZN(
        n14319) );
  AOI221_X2 U6660 ( .B1(n17526), .B2(n25870), .C1(n25867), .C2(n25469), .A(
        n14344), .ZN(n14342) );
  AOI221_X2 U6663 ( .B1(n25859), .B2(n25649), .C1(n25857), .C2(n25162), .A(
        n14350), .ZN(n14341) );
  OAI22_X2 U6664 ( .A1(n17557), .A2(n25855), .B1(n17529), .B2(n25853), .ZN(
        n14350) );
  AOI221_X2 U6667 ( .B1(n17549), .B2(n25852), .C1(n17540), .C2(n25849), .A(
        n14351), .ZN(n14340) );
  AOI221_X2 U6669 ( .B1(n17550), .B2(n25842), .C1(n17541), .C2(n25839), .A(
        n14352), .ZN(n14339) );
  OAI22_X2 U6670 ( .A1(n25838), .A2(n27095), .B1(n25835), .B2(n27159), .ZN(
        n14352) );
  NAND4_X2 U6673 ( .A1(n14358), .A2(n14359), .A3(n14360), .A4(n14361), .ZN(
        n14357) );
  AOI221_X2 U6674 ( .B1(n25906), .B2(n25002), .C1(n25903), .C2(n25468), .A(
        n14364), .ZN(n14361) );
  AOI221_X2 U6678 ( .B1(n25896), .B2(n25001), .C1(n25893), .C2(n25467), .A(
        n14369), .ZN(n14360) );
  OAI22_X2 U6679 ( .A1(n17515), .A2(n25891), .B1(n17487), .B2(n25889), .ZN(
        n14369) );
  AOI221_X2 U6682 ( .B1(n17500), .B2(n25888), .C1(n17491), .C2(n25886), .A(
        n14370), .ZN(n14359) );
  AOI221_X2 U6684 ( .B1(n17517), .B2(n25878), .C1(n17508), .C2(n25875), .A(
        n14373), .ZN(n14358) );
  OAI22_X2 U6685 ( .A1(n25874), .A2(n26520), .B1(n25871), .B2(n26616), .ZN(
        n14373) );
  NAND4_X2 U6686 ( .A1(n14376), .A2(n14377), .A3(n14378), .A4(n14379), .ZN(
        n14356) );
  AOI221_X2 U6687 ( .B1(n17489), .B2(n25870), .C1(n25867), .C2(n25466), .A(
        n14381), .ZN(n14379) );
  AOI221_X2 U6690 ( .B1(n25860), .B2(n25648), .C1(n25857), .C2(n25161), .A(
        n14387), .ZN(n14378) );
  OAI22_X2 U6691 ( .A1(n17520), .A2(n25856), .B1(n17492), .B2(n25853), .ZN(
        n14387) );
  AOI221_X2 U6694 ( .B1(n17512), .B2(n25852), .C1(n17503), .C2(n25849), .A(
        n14388), .ZN(n14377) );
  AOI221_X2 U6696 ( .B1(n17513), .B2(n25842), .C1(n17504), .C2(n25839), .A(
        n14389), .ZN(n14376) );
  OAI22_X2 U6697 ( .A1(n25838), .A2(n27096), .B1(n25836), .B2(n27160), .ZN(
        n14389) );
  NAND4_X2 U6700 ( .A1(n14395), .A2(n14396), .A3(n14397), .A4(n14398), .ZN(
        n14394) );
  AOI221_X2 U6701 ( .B1(n25905), .B2(n25000), .C1(n25903), .C2(n25465), .A(
        n14401), .ZN(n14398) );
  AOI221_X2 U6705 ( .B1(n25896), .B2(n24999), .C1(n25893), .C2(n25464), .A(
        n14406), .ZN(n14397) );
  OAI22_X2 U6706 ( .A1(n17478), .A2(n25891), .B1(n17450), .B2(n25889), .ZN(
        n14406) );
  AOI221_X2 U6709 ( .B1(n17463), .B2(n25888), .C1(n17454), .C2(n25886), .A(
        n14407), .ZN(n14396) );
  AOI221_X2 U6711 ( .B1(n17480), .B2(n25878), .C1(n17471), .C2(n25875), .A(
        n14410), .ZN(n14395) );
  OAI22_X2 U6712 ( .A1(n25874), .A2(n26521), .B1(n25871), .B2(n26617), .ZN(
        n14410) );
  NAND4_X2 U6713 ( .A1(n14413), .A2(n14414), .A3(n14415), .A4(n14416), .ZN(
        n14393) );
  AOI221_X2 U6714 ( .B1(n17452), .B2(n25870), .C1(n25867), .C2(n25463), .A(
        n14418), .ZN(n14416) );
  AOI221_X2 U6717 ( .B1(n25859), .B2(n25647), .C1(n25857), .C2(n25160), .A(
        n14424), .ZN(n14415) );
  OAI22_X2 U6718 ( .A1(n17483), .A2(n25856), .B1(n17455), .B2(n25853), .ZN(
        n14424) );
  AOI221_X2 U6721 ( .B1(n17475), .B2(n25852), .C1(n17466), .C2(n25849), .A(
        n14425), .ZN(n14414) );
  AOI221_X2 U6723 ( .B1(n17476), .B2(n25842), .C1(n17467), .C2(n25839), .A(
        n14426), .ZN(n14413) );
  OAI22_X2 U6724 ( .A1(n25838), .A2(n27097), .B1(n25835), .B2(n27161), .ZN(
        n14426) );
  NAND4_X2 U6727 ( .A1(n14432), .A2(n14433), .A3(n14434), .A4(n14435), .ZN(
        n14431) );
  AOI221_X2 U6728 ( .B1(n25906), .B2(n24998), .C1(n25903), .C2(n25462), .A(
        n14438), .ZN(n14435) );
  AOI221_X2 U6732 ( .B1(n25896), .B2(n24997), .C1(n25893), .C2(n25461), .A(
        n14443), .ZN(n14434) );
  OAI22_X2 U6733 ( .A1(n17441), .A2(n25891), .B1(n17413), .B2(n25889), .ZN(
        n14443) );
  AOI221_X2 U6736 ( .B1(n17426), .B2(n25888), .C1(n17417), .C2(n25886), .A(
        n14444), .ZN(n14433) );
  AOI221_X2 U6738 ( .B1(n17443), .B2(n25878), .C1(n17434), .C2(n25875), .A(
        n14447), .ZN(n14432) );
  OAI22_X2 U6739 ( .A1(n25874), .A2(n26522), .B1(n25871), .B2(n26618), .ZN(
        n14447) );
  NAND4_X2 U6740 ( .A1(n14450), .A2(n14451), .A3(n14452), .A4(n14453), .ZN(
        n14430) );
  AOI221_X2 U6741 ( .B1(n17415), .B2(n25870), .C1(n25867), .C2(n25460), .A(
        n14455), .ZN(n14453) );
  AOI221_X2 U6744 ( .B1(n25860), .B2(n25646), .C1(n25857), .C2(n25159), .A(
        n14461), .ZN(n14452) );
  OAI22_X2 U6745 ( .A1(n17446), .A2(n25855), .B1(n17418), .B2(n25853), .ZN(
        n14461) );
  AOI221_X2 U6748 ( .B1(n17438), .B2(n25852), .C1(n17429), .C2(n25849), .A(
        n14462), .ZN(n14451) );
  AOI221_X2 U6750 ( .B1(n17439), .B2(n25842), .C1(n17430), .C2(n25839), .A(
        n14463), .ZN(n14450) );
  OAI22_X2 U6751 ( .A1(n25838), .A2(n27098), .B1(n25835), .B2(n27162), .ZN(
        n14463) );
  NAND4_X2 U6754 ( .A1(n14469), .A2(n14470), .A3(n14471), .A4(n14472), .ZN(
        n14468) );
  AOI221_X2 U6755 ( .B1(n25905), .B2(n24996), .C1(n25903), .C2(n25459), .A(
        n14475), .ZN(n14472) );
  AOI221_X2 U6759 ( .B1(n25896), .B2(n24995), .C1(n25893), .C2(n25458), .A(
        n14480), .ZN(n14471) );
  OAI22_X2 U6760 ( .A1(n17404), .A2(n25891), .B1(n17376), .B2(n25890), .ZN(
        n14480) );
  AOI221_X2 U6763 ( .B1(n17389), .B2(n25888), .C1(n17380), .C2(n25886), .A(
        n14481), .ZN(n14470) );
  AOI221_X2 U6765 ( .B1(n17406), .B2(n25878), .C1(n17397), .C2(n25875), .A(
        n14484), .ZN(n14469) );
  OAI22_X2 U6766 ( .A1(n25874), .A2(n26523), .B1(n25872), .B2(n26619), .ZN(
        n14484) );
  NAND4_X2 U6767 ( .A1(n14487), .A2(n14488), .A3(n14489), .A4(n14490), .ZN(
        n14467) );
  AOI221_X2 U6768 ( .B1(n17378), .B2(n25870), .C1(n25867), .C2(n25457), .A(
        n14492), .ZN(n14490) );
  AOI221_X2 U6771 ( .B1(n25859), .B2(n25645), .C1(n25857), .C2(n25158), .A(
        n14498), .ZN(n14489) );
  OAI22_X2 U6772 ( .A1(n17409), .A2(n25855), .B1(n17381), .B2(n25854), .ZN(
        n14498) );
  AOI221_X2 U6775 ( .B1(n17401), .B2(n25852), .C1(n17392), .C2(n25849), .A(
        n14499), .ZN(n14488) );
  AOI221_X2 U6777 ( .B1(n17402), .B2(n25842), .C1(n17393), .C2(n25839), .A(
        n14500), .ZN(n14487) );
  OAI22_X2 U6778 ( .A1(n25837), .A2(n27099), .B1(n25836), .B2(n27163), .ZN(
        n14500) );
  NAND4_X2 U6781 ( .A1(n14506), .A2(n14507), .A3(n14508), .A4(n14509), .ZN(
        n14505) );
  AOI221_X2 U6782 ( .B1(n25906), .B2(n24994), .C1(n25903), .C2(n25456), .A(
        n14512), .ZN(n14509) );
  AOI221_X2 U6786 ( .B1(n25896), .B2(n24993), .C1(n25893), .C2(n25455), .A(
        n14517), .ZN(n14508) );
  OAI22_X2 U6787 ( .A1(n17367), .A2(n25892), .B1(n17339), .B2(n25890), .ZN(
        n14517) );
  AOI221_X2 U6790 ( .B1(n17352), .B2(n25888), .C1(n17343), .C2(n25886), .A(
        n14518), .ZN(n14507) );
  AOI221_X2 U6792 ( .B1(n17369), .B2(n25878), .C1(n17360), .C2(n25875), .A(
        n14521), .ZN(n14506) );
  OAI22_X2 U6793 ( .A1(n25874), .A2(n26524), .B1(n25872), .B2(n26620), .ZN(
        n14521) );
  NAND4_X2 U6794 ( .A1(n14524), .A2(n14525), .A3(n14526), .A4(n14527), .ZN(
        n14504) );
  AOI221_X2 U6795 ( .B1(n17341), .B2(n25870), .C1(n25867), .C2(n25454), .A(
        n14529), .ZN(n14527) );
  AOI221_X2 U6798 ( .B1(n25860), .B2(n25644), .C1(n25857), .C2(n25157), .A(
        n14535), .ZN(n14526) );
  OAI22_X2 U6799 ( .A1(n17372), .A2(n25856), .B1(n17344), .B2(n25854), .ZN(
        n14535) );
  AOI221_X2 U6802 ( .B1(n17364), .B2(n25852), .C1(n17355), .C2(n25849), .A(
        n14536), .ZN(n14525) );
  AOI221_X2 U6804 ( .B1(n17365), .B2(n25842), .C1(n17356), .C2(n25839), .A(
        n14537), .ZN(n14524) );
  OAI22_X2 U6805 ( .A1(n25838), .A2(n27100), .B1(n25836), .B2(n27164), .ZN(
        n14537) );
  NAND4_X2 U6808 ( .A1(n14543), .A2(n14544), .A3(n14545), .A4(n14546), .ZN(
        n14542) );
  AOI221_X2 U6809 ( .B1(n25905), .B2(n24992), .C1(n25903), .C2(n25453), .A(
        n14549), .ZN(n14546) );
  AOI221_X2 U6813 ( .B1(n25896), .B2(n24991), .C1(n25893), .C2(n25452), .A(
        n14554), .ZN(n14545) );
  OAI22_X2 U6814 ( .A1(n17330), .A2(n25891), .B1(n17302), .B2(n25890), .ZN(
        n14554) );
  AOI221_X2 U6817 ( .B1(n17315), .B2(n25888), .C1(n17306), .C2(n25886), .A(
        n14555), .ZN(n14544) );
  AOI221_X2 U6819 ( .B1(n17332), .B2(n25878), .C1(n17323), .C2(n25875), .A(
        n14558), .ZN(n14543) );
  OAI22_X2 U6820 ( .A1(n25874), .A2(n26525), .B1(n25872), .B2(n26621), .ZN(
        n14558) );
  NAND4_X2 U6821 ( .A1(n14561), .A2(n14562), .A3(n14563), .A4(n14564), .ZN(
        n14541) );
  AOI221_X2 U6822 ( .B1(n17304), .B2(n25870), .C1(n25867), .C2(n25451), .A(
        n14566), .ZN(n14564) );
  AOI221_X2 U6825 ( .B1(n25860), .B2(n25643), .C1(n25857), .C2(n25156), .A(
        n14572), .ZN(n14563) );
  OAI22_X2 U6826 ( .A1(n17335), .A2(n25855), .B1(n17307), .B2(n25854), .ZN(
        n14572) );
  AOI221_X2 U6829 ( .B1(n17327), .B2(n25852), .C1(n17318), .C2(n25849), .A(
        n14573), .ZN(n14562) );
  AOI221_X2 U6831 ( .B1(n17328), .B2(n25842), .C1(n17319), .C2(n25839), .A(
        n14574), .ZN(n14561) );
  OAI22_X2 U6832 ( .A1(n25837), .A2(n27101), .B1(n25836), .B2(n27165), .ZN(
        n14574) );
  NAND4_X2 U6835 ( .A1(n14580), .A2(n14581), .A3(n14582), .A4(n14583), .ZN(
        n14579) );
  AOI221_X2 U6836 ( .B1(n25906), .B2(n24990), .C1(n25903), .C2(n25450), .A(
        n14586), .ZN(n14583) );
  AOI221_X2 U6840 ( .B1(n25895), .B2(n24989), .C1(n25893), .C2(n25449), .A(
        n14591), .ZN(n14582) );
  OAI22_X2 U6841 ( .A1(n17293), .A2(n25892), .B1(n17265), .B2(n25890), .ZN(
        n14591) );
  AOI221_X2 U6844 ( .B1(n17278), .B2(n25887), .C1(n17269), .C2(n25885), .A(
        n14592), .ZN(n14581) );
  AOI221_X2 U6846 ( .B1(n17295), .B2(n25877), .C1(n17286), .C2(n25875), .A(
        n14595), .ZN(n14580) );
  OAI22_X2 U6847 ( .A1(n25874), .A2(n26526), .B1(n25872), .B2(n26622), .ZN(
        n14595) );
  NAND4_X2 U6848 ( .A1(n14598), .A2(n14599), .A3(n14600), .A4(n14601), .ZN(
        n14578) );
  AOI221_X2 U6849 ( .B1(n17267), .B2(n25870), .C1(n25867), .C2(n25448), .A(
        n14603), .ZN(n14601) );
  AOI221_X2 U6852 ( .B1(n25860), .B2(n25642), .C1(n25857), .C2(n25155), .A(
        n14609), .ZN(n14600) );
  OAI22_X2 U6853 ( .A1(n17298), .A2(n25856), .B1(n17270), .B2(n25854), .ZN(
        n14609) );
  AOI221_X2 U6856 ( .B1(n17290), .B2(n25851), .C1(n17281), .C2(n25849), .A(
        n14610), .ZN(n14599) );
  AOI221_X2 U6858 ( .B1(n17291), .B2(n25841), .C1(n17282), .C2(n25839), .A(
        n14611), .ZN(n14598) );
  OAI22_X2 U6859 ( .A1(n25838), .A2(n27102), .B1(n25836), .B2(n27166), .ZN(
        n14611) );
  NAND4_X2 U6862 ( .A1(n14617), .A2(n14618), .A3(n14619), .A4(n14620), .ZN(
        n14616) );
  AOI221_X2 U6863 ( .B1(n25906), .B2(n24988), .C1(n25904), .C2(n25447), .A(
        n14623), .ZN(n14620) );
  AOI221_X2 U6867 ( .B1(n25896), .B2(n24987), .C1(n25893), .C2(n25446), .A(
        n14628), .ZN(n14619) );
  OAI22_X2 U6868 ( .A1(n17256), .A2(n25892), .B1(n17228), .B2(n25890), .ZN(
        n14628) );
  AOI221_X2 U6871 ( .B1(n17241), .B2(n25888), .C1(n17232), .C2(n25886), .A(
        n14629), .ZN(n14618) );
  AOI221_X2 U6873 ( .B1(n17258), .B2(n25878), .C1(n17249), .C2(n25876), .A(
        n14632), .ZN(n14617) );
  OAI22_X2 U6874 ( .A1(n25874), .A2(n26527), .B1(n25872), .B2(n26623), .ZN(
        n14632) );
  NAND4_X2 U6875 ( .A1(n14635), .A2(n14636), .A3(n14637), .A4(n14638), .ZN(
        n14615) );
  AOI221_X2 U6876 ( .B1(n17230), .B2(n25869), .C1(n25868), .C2(n25445), .A(
        n14640), .ZN(n14638) );
  AOI221_X2 U6879 ( .B1(n25860), .B2(n25641), .C1(n25858), .C2(n25154), .A(
        n14646), .ZN(n14637) );
  OAI22_X2 U6880 ( .A1(n17261), .A2(n25855), .B1(n17233), .B2(n25854), .ZN(
        n14646) );
  AOI221_X2 U6883 ( .B1(n17253), .B2(n25852), .C1(n17244), .C2(n25850), .A(
        n14647), .ZN(n14636) );
  AOI221_X2 U6885 ( .B1(n17254), .B2(n25842), .C1(n17245), .C2(n25840), .A(
        n14648), .ZN(n14635) );
  OAI22_X2 U6886 ( .A1(n25837), .A2(n27103), .B1(n25836), .B2(n27167), .ZN(
        n14648) );
  NAND4_X2 U6889 ( .A1(n14654), .A2(n14655), .A3(n14656), .A4(n14657), .ZN(
        n14653) );
  AOI221_X2 U6890 ( .B1(n25905), .B2(n24986), .C1(n25903), .C2(n25444), .A(
        n14660), .ZN(n14657) );
  AOI221_X2 U6894 ( .B1(n25895), .B2(n24985), .C1(n25894), .C2(n25443), .A(
        n14665), .ZN(n14656) );
  OAI22_X2 U6895 ( .A1(n17219), .A2(n25891), .B1(n17191), .B2(n25890), .ZN(
        n14665) );
  AOI221_X2 U6898 ( .B1(n17204), .B2(n25887), .C1(n17195), .C2(n25885), .A(
        n14666), .ZN(n14655) );
  AOI221_X2 U6900 ( .B1(n17221), .B2(n25877), .C1(n17212), .C2(n25876), .A(
        n14669), .ZN(n14654) );
  OAI22_X2 U6901 ( .A1(n25874), .A2(n26528), .B1(n25872), .B2(n26624), .ZN(
        n14669) );
  NAND4_X2 U6902 ( .A1(n14672), .A2(n14673), .A3(n14674), .A4(n14675), .ZN(
        n14652) );
  AOI221_X2 U6903 ( .B1(n17193), .B2(n25870), .C1(n25867), .C2(n25442), .A(
        n14677), .ZN(n14675) );
  AOI221_X2 U6906 ( .B1(n25859), .B2(n25640), .C1(n25857), .C2(n25153), .A(
        n14683), .ZN(n14674) );
  OAI22_X2 U6907 ( .A1(n17224), .A2(n25855), .B1(n17196), .B2(n25854), .ZN(
        n14683) );
  AOI221_X2 U6910 ( .B1(n17216), .B2(n25851), .C1(n17207), .C2(n25849), .A(
        n14684), .ZN(n14673) );
  AOI221_X2 U6912 ( .B1(n17217), .B2(n25841), .C1(n17208), .C2(n25840), .A(
        n14685), .ZN(n14672) );
  OAI22_X2 U6913 ( .A1(n25838), .A2(n27104), .B1(n25836), .B2(n27168), .ZN(
        n14685) );
  NAND4_X2 U6916 ( .A1(n14691), .A2(n14692), .A3(n14693), .A4(n14694), .ZN(
        n14690) );
  AOI221_X2 U6917 ( .B1(n25905), .B2(n24984), .C1(n25904), .C2(n25441), .A(
        n14697), .ZN(n14694) );
  AOI221_X2 U6921 ( .B1(n25896), .B2(n24983), .C1(n25894), .C2(n25440), .A(
        n14702), .ZN(n14693) );
  OAI22_X2 U6922 ( .A1(n17182), .A2(n25892), .B1(n17154), .B2(n25890), .ZN(
        n14702) );
  AOI221_X2 U6925 ( .B1(n17167), .B2(n25887), .C1(n17158), .C2(n25886), .A(
        n14703), .ZN(n14692) );
  AOI221_X2 U6927 ( .B1(n17184), .B2(n25878), .C1(n17175), .C2(n25875), .A(
        n14706), .ZN(n14691) );
  OAI22_X2 U6928 ( .A1(n25874), .A2(n26529), .B1(n25872), .B2(n26625), .ZN(
        n14706) );
  NAND4_X2 U6929 ( .A1(n14709), .A2(n14710), .A3(n14711), .A4(n14712), .ZN(
        n14689) );
  AOI221_X2 U6930 ( .B1(n17156), .B2(n25869), .C1(n25868), .C2(n25439), .A(
        n14714), .ZN(n14712) );
  AOI221_X2 U6933 ( .B1(n25859), .B2(n25639), .C1(n25858), .C2(n25152), .A(
        n14720), .ZN(n14711) );
  OAI22_X2 U6934 ( .A1(n17187), .A2(n25856), .B1(n17159), .B2(n25854), .ZN(
        n14720) );
  AOI221_X2 U6937 ( .B1(n17179), .B2(n25852), .C1(n17170), .C2(n25850), .A(
        n14721), .ZN(n14710) );
  AOI221_X2 U6939 ( .B1(n17180), .B2(n25842), .C1(n17171), .C2(n25839), .A(
        n14722), .ZN(n14709) );
  OAI22_X2 U6940 ( .A1(n25837), .A2(n27105), .B1(n25836), .B2(n27169), .ZN(
        n14722) );
  NAND4_X2 U6943 ( .A1(n14728), .A2(n14729), .A3(n14730), .A4(n14731), .ZN(
        n14727) );
  AOI221_X2 U6944 ( .B1(n25906), .B2(n24982), .C1(n25903), .C2(n25438), .A(
        n14734), .ZN(n14731) );
  AOI221_X2 U6948 ( .B1(n25896), .B2(n24981), .C1(n25893), .C2(n25437), .A(
        n14739), .ZN(n14730) );
  OAI22_X2 U6949 ( .A1(n17145), .A2(n25891), .B1(n17117), .B2(n25890), .ZN(
        n14739) );
  AOI221_X2 U6952 ( .B1(n17130), .B2(n25887), .C1(n17121), .C2(n25885), .A(
        n14740), .ZN(n14729) );
  AOI221_X2 U6954 ( .B1(n17147), .B2(n25878), .C1(n17138), .C2(n25876), .A(
        n14743), .ZN(n14728) );
  OAI22_X2 U6955 ( .A1(n25874), .A2(n26530), .B1(n25872), .B2(n26626), .ZN(
        n14743) );
  NAND4_X2 U6956 ( .A1(n14746), .A2(n14747), .A3(n14748), .A4(n14749), .ZN(
        n14726) );
  AOI221_X2 U6957 ( .B1(n17119), .B2(n25869), .C1(n25867), .C2(n25436), .A(
        n14751), .ZN(n14749) );
  AOI221_X2 U6960 ( .B1(n25860), .B2(n25638), .C1(n25857), .C2(n25151), .A(
        n14757), .ZN(n14748) );
  OAI22_X2 U6961 ( .A1(n17150), .A2(n25856), .B1(n17122), .B2(n25854), .ZN(
        n14757) );
  AOI221_X2 U6964 ( .B1(n17142), .B2(n25852), .C1(n17133), .C2(n25849), .A(
        n14758), .ZN(n14747) );
  AOI221_X2 U6966 ( .B1(n17143), .B2(n25842), .C1(n17134), .C2(n25840), .A(
        n14759), .ZN(n14746) );
  OAI22_X2 U6967 ( .A1(n25838), .A2(n27106), .B1(n25836), .B2(n27170), .ZN(
        n14759) );
  OAI22_X2 U6968 ( .A1(n17114), .A2(n25907), .B1(n14762), .B2(n12153), .ZN(
        n23496) );
  NOR2_X2 U6969 ( .A1(n14763), .A2(n14764), .ZN(n14762) );
  NAND4_X2 U6970 ( .A1(n14765), .A2(n14766), .A3(n14767), .A4(n14768), .ZN(
        n14764) );
  AOI221_X2 U6971 ( .B1(n25906), .B2(n25637), .C1(n25903), .C2(n25150), .A(
        n14771), .ZN(n14768) );
  AOI221_X2 U6975 ( .B1(n25896), .B2(n25636), .C1(n25893), .C2(n25149), .A(
        n14776), .ZN(n14767) );
  OAI22_X2 U6976 ( .A1(n17108), .A2(n25891), .B1(n17080), .B2(n25890), .ZN(
        n14776) );
  AOI221_X2 U6979 ( .B1(n17093), .B2(n25887), .C1(n17084), .C2(n25885), .A(
        n14777), .ZN(n14766) );
  AOI221_X2 U6981 ( .B1(n17110), .B2(n25878), .C1(n17101), .C2(n25876), .A(
        n14780), .ZN(n14765) );
  OAI22_X2 U6982 ( .A1(n25874), .A2(n26531), .B1(n25872), .B2(n26627), .ZN(
        n14780) );
  NAND4_X2 U6983 ( .A1(n14783), .A2(n14784), .A3(n14785), .A4(n14786), .ZN(
        n14763) );
  AOI221_X2 U6984 ( .B1(n17082), .B2(n25869), .C1(n25867), .C2(n25435), .A(
        n14788), .ZN(n14786) );
  AOI221_X2 U6987 ( .B1(n25860), .B2(n25635), .C1(n25858), .C2(n25148), .A(
        n14794), .ZN(n14785) );
  OAI22_X2 U6988 ( .A1(n17113), .A2(n25855), .B1(n17085), .B2(n25854), .ZN(
        n14794) );
  AOI221_X2 U6991 ( .B1(n17105), .B2(n25852), .C1(n17096), .C2(n25850), .A(
        n14795), .ZN(n14784) );
  AOI221_X2 U6993 ( .B1(n17106), .B2(n25842), .C1(n17097), .C2(n25840), .A(
        n14796), .ZN(n14783) );
  OAI22_X2 U6994 ( .A1(n25838), .A2(n27107), .B1(n25836), .B2(n27171), .ZN(
        n14796) );
  OAI22_X2 U6995 ( .A1(n17077), .A2(n25909), .B1(n14799), .B2(n12153), .ZN(
        n23497) );
  NOR2_X2 U6996 ( .A1(n14800), .A2(n14801), .ZN(n14799) );
  NAND4_X2 U6997 ( .A1(n14802), .A2(n14803), .A3(n14804), .A4(n14805), .ZN(
        n14801) );
  AOI221_X2 U6998 ( .B1(n25906), .B2(n25634), .C1(n25904), .C2(n25147), .A(
        n14808), .ZN(n14805) );
  AOI221_X2 U7002 ( .B1(n25896), .B2(n25633), .C1(n25894), .C2(n25146), .A(
        n14813), .ZN(n14804) );
  OAI22_X2 U7003 ( .A1(n17071), .A2(n25891), .B1(n17043), .B2(n25890), .ZN(
        n14813) );
  AOI221_X2 U7006 ( .B1(n17056), .B2(n25888), .C1(n17047), .C2(n25885), .A(
        n14814), .ZN(n14803) );
  AOI221_X2 U7008 ( .B1(n17073), .B2(n25878), .C1(n17064), .C2(n25875), .A(
        n14817), .ZN(n14802) );
  OAI22_X2 U7009 ( .A1(n25874), .A2(n26532), .B1(n25872), .B2(n26628), .ZN(
        n14817) );
  NAND4_X2 U7010 ( .A1(n14820), .A2(n14821), .A3(n14822), .A4(n14823), .ZN(
        n14800) );
  AOI221_X2 U7011 ( .B1(n17045), .B2(n25869), .C1(n25868), .C2(n25434), .A(
        n14825), .ZN(n14823) );
  AOI221_X2 U7014 ( .B1(n25860), .B2(n25632), .C1(n25857), .C2(n25145), .A(
        n14831), .ZN(n14822) );
  OAI22_X2 U7015 ( .A1(n17076), .A2(n25855), .B1(n17048), .B2(n25854), .ZN(
        n14831) );
  AOI221_X2 U7018 ( .B1(n17068), .B2(n25852), .C1(n17059), .C2(n25849), .A(
        n14832), .ZN(n14821) );
  AOI221_X2 U7020 ( .B1(n17069), .B2(n25842), .C1(n17060), .C2(n25839), .A(
        n14833), .ZN(n14820) );
  OAI22_X2 U7021 ( .A1(n25838), .A2(n27108), .B1(n25836), .B2(n27172), .ZN(
        n14833) );
  OAI22_X2 U7022 ( .A1(n17040), .A2(n25907), .B1(n14836), .B2(n12153), .ZN(
        n23498) );
  NOR2_X2 U7023 ( .A1(n14837), .A2(n14838), .ZN(n14836) );
  NAND4_X2 U7024 ( .A1(n14839), .A2(n14840), .A3(n14841), .A4(n14842), .ZN(
        n14838) );
  AOI221_X2 U7025 ( .B1(n25905), .B2(n25631), .C1(n25904), .C2(n25144), .A(
        n14845), .ZN(n14842) );
  AOI221_X2 U7029 ( .B1(n25895), .B2(n25630), .C1(n25894), .C2(n25143), .A(
        n14850), .ZN(n14841) );
  OAI22_X2 U7030 ( .A1(n17034), .A2(n25892), .B1(n17006), .B2(n25890), .ZN(
        n14850) );
  AOI221_X2 U7033 ( .B1(n17019), .B2(n25888), .C1(n17010), .C2(n25886), .A(
        n14851), .ZN(n14840) );
  AOI221_X2 U7035 ( .B1(n17036), .B2(n25877), .C1(n17027), .C2(n25875), .A(
        n14854), .ZN(n14839) );
  OAI22_X2 U7036 ( .A1(n25874), .A2(n26533), .B1(n25872), .B2(n26629), .ZN(
        n14854) );
  NAND4_X2 U7037 ( .A1(n14857), .A2(n14858), .A3(n14859), .A4(n14860), .ZN(
        n14837) );
  AOI221_X2 U7038 ( .B1(n17008), .B2(n25870), .C1(n25867), .C2(n25433), .A(
        n14862), .ZN(n14860) );
  AOI221_X2 U7041 ( .B1(n25859), .B2(n25629), .C1(n25857), .C2(n25142), .A(
        n14868), .ZN(n14859) );
  OAI22_X2 U7042 ( .A1(n17039), .A2(n25856), .B1(n17011), .B2(n25854), .ZN(
        n14868) );
  AOI221_X2 U7045 ( .B1(n17031), .B2(n25851), .C1(n17022), .C2(n25849), .A(
        n14869), .ZN(n14858) );
  AOI221_X2 U7047 ( .B1(n17032), .B2(n25841), .C1(n17023), .C2(n25839), .A(
        n14870), .ZN(n14857) );
  OAI22_X2 U7048 ( .A1(n25837), .A2(n27109), .B1(n25836), .B2(n27173), .ZN(
        n14870) );
  OAI22_X2 U7049 ( .A1(n17003), .A2(n25907), .B1(n14873), .B2(n12153), .ZN(
        n23499) );
  NOR2_X2 U7050 ( .A1(n14874), .A2(n14875), .ZN(n14873) );
  NAND4_X2 U7051 ( .A1(n14876), .A2(n14877), .A3(n14878), .A4(n14879), .ZN(
        n14875) );
  AOI221_X2 U7052 ( .B1(n25905), .B2(n25628), .C1(n25903), .C2(n25141), .A(
        n14882), .ZN(n14879) );
  AOI221_X2 U7056 ( .B1(n25895), .B2(n25627), .C1(n25893), .C2(n25140), .A(
        n14887), .ZN(n14878) );
  OAI22_X2 U7057 ( .A1(n16997), .A2(n25891), .B1(n16969), .B2(n25890), .ZN(
        n14887) );
  AOI221_X2 U7060 ( .B1(n16982), .B2(n25887), .C1(n16973), .C2(n25886), .A(
        n14888), .ZN(n14877) );
  AOI221_X2 U7062 ( .B1(n16999), .B2(n25877), .C1(n16990), .C2(n25876), .A(
        n14891), .ZN(n14876) );
  OAI22_X2 U7063 ( .A1(n25874), .A2(n26534), .B1(n25872), .B2(n26630), .ZN(
        n14891) );
  NAND4_X2 U7064 ( .A1(n14894), .A2(n14895), .A3(n14896), .A4(n14897), .ZN(
        n14874) );
  AOI221_X2 U7065 ( .B1(n16971), .B2(n25870), .C1(n25868), .C2(n25432), .A(
        n14899), .ZN(n14897) );
  AOI221_X2 U7068 ( .B1(n25859), .B2(n25626), .C1(n25858), .C2(n25139), .A(
        n14905), .ZN(n14896) );
  OAI22_X2 U7069 ( .A1(n17002), .A2(n25855), .B1(n16974), .B2(n25854), .ZN(
        n14905) );
  AOI221_X2 U7072 ( .B1(n16994), .B2(n25851), .C1(n16985), .C2(n25849), .A(
        n14906), .ZN(n14895) );
  AOI221_X2 U7074 ( .B1(n16995), .B2(n25841), .C1(n16986), .C2(n25840), .A(
        n14907), .ZN(n14894) );
  OAI22_X2 U7075 ( .A1(n25837), .A2(n27110), .B1(n25836), .B2(n27174), .ZN(
        n14907) );
  NAND4_X2 U7078 ( .A1(n14913), .A2(n14914), .A3(n14915), .A4(n14916), .ZN(
        n14912) );
  AOI221_X2 U7079 ( .B1(n25906), .B2(n24980), .C1(n25903), .C2(n25431), .A(
        n14919), .ZN(n14916) );
  AOI221_X2 U7083 ( .B1(n25896), .B2(n24979), .C1(n25894), .C2(n25430), .A(
        n14924), .ZN(n14915) );
  OAI22_X2 U7084 ( .A1(n16960), .A2(n25892), .B1(n16932), .B2(n25889), .ZN(
        n14924) );
  AOI221_X2 U7087 ( .B1(n16945), .B2(n25887), .C1(n16936), .C2(n25886), .A(
        n14925), .ZN(n14914) );
  AOI221_X2 U7089 ( .B1(n16962), .B2(n25878), .C1(n16953), .C2(n25875), .A(
        n14928), .ZN(n14913) );
  OAI22_X2 U7090 ( .A1(n25874), .A2(n26535), .B1(n25871), .B2(n26631), .ZN(
        n14928) );
  NAND4_X2 U7091 ( .A1(n14931), .A2(n14932), .A3(n14933), .A4(n14934), .ZN(
        n14911) );
  AOI221_X2 U7092 ( .B1(n16934), .B2(n25869), .C1(n25868), .C2(n25429), .A(
        n14936), .ZN(n14934) );
  AOI221_X2 U7095 ( .B1(n25860), .B2(n25625), .C1(n25858), .C2(n25138), .A(
        n14942), .ZN(n14933) );
  OAI22_X2 U7096 ( .A1(n16965), .A2(n25856), .B1(n16937), .B2(n25853), .ZN(
        n14942) );
  AOI221_X2 U7099 ( .B1(n16957), .B2(n25852), .C1(n16948), .C2(n25849), .A(
        n14943), .ZN(n14932) );
  AOI221_X2 U7101 ( .B1(n16958), .B2(n25842), .C1(n16949), .C2(n25839), .A(
        n14944), .ZN(n14931) );
  OAI22_X2 U7102 ( .A1(n25837), .A2(n27143), .B1(n25835), .B2(n27207), .ZN(
        n14944) );
  NAND4_X2 U7105 ( .A1(n14950), .A2(n14951), .A3(n14952), .A4(n14953), .ZN(
        n14949) );
  AOI221_X2 U7106 ( .B1(n25905), .B2(n24978), .C1(n25903), .C2(n25428), .A(
        n14956), .ZN(n14953) );
  AOI221_X2 U7110 ( .B1(n25895), .B2(n24977), .C1(n25893), .C2(n25427), .A(
        n14961), .ZN(n14952) );
  OAI22_X2 U7111 ( .A1(n16923), .A2(n25892), .B1(n16895), .B2(n25890), .ZN(
        n14961) );
  AOI221_X2 U7114 ( .B1(n16908), .B2(n25887), .C1(n16899), .C2(n25885), .A(
        n14962), .ZN(n14951) );
  AOI221_X2 U7116 ( .B1(n16925), .B2(n25877), .C1(n16916), .C2(n25875), .A(
        n14965), .ZN(n14950) );
  OAI22_X2 U7117 ( .A1(n25874), .A2(n26536), .B1(n25872), .B2(n26632), .ZN(
        n14965) );
  NAND4_X2 U7118 ( .A1(n14968), .A2(n14969), .A3(n14970), .A4(n14971), .ZN(
        n14948) );
  AOI221_X2 U7119 ( .B1(n16897), .B2(n25870), .C1(n25867), .C2(n25426), .A(
        n14973), .ZN(n14971) );
  AOI221_X2 U7122 ( .B1(n25859), .B2(n24976), .C1(n25857), .C2(n25425), .A(
        n14979), .ZN(n14970) );
  OAI22_X2 U7123 ( .A1(n16928), .A2(n25855), .B1(n16900), .B2(n25854), .ZN(
        n14979) );
  AOI221_X2 U7126 ( .B1(n16920), .B2(n25851), .C1(n16911), .C2(n25849), .A(
        n14980), .ZN(n14969) );
  AOI221_X2 U7128 ( .B1(n16921), .B2(n25841), .C1(n16912), .C2(n25839), .A(
        n14981), .ZN(n14968) );
  OAI22_X2 U7129 ( .A1(n25837), .A2(n27144), .B1(n25836), .B2(n27208), .ZN(
        n14981) );
  NAND4_X2 U7132 ( .A1(n14987), .A2(n14988), .A3(n14989), .A4(n14990), .ZN(
        n14986) );
  AOI221_X2 U7133 ( .B1(n25905), .B2(n24975), .C1(n25904), .C2(n25424), .A(
        n14993), .ZN(n14990) );
  AOI221_X2 U7137 ( .B1(n25896), .B2(n24974), .C1(n25893), .C2(n25423), .A(
        n14998), .ZN(n14989) );
  OAI22_X2 U7138 ( .A1(n16886), .A2(n25892), .B1(n16858), .B2(n25889), .ZN(
        n14998) );
  AOI221_X2 U7141 ( .B1(n16871), .B2(n25887), .C1(n16862), .C2(n25885), .A(
        n14999), .ZN(n14988) );
  AOI221_X2 U7143 ( .B1(n16888), .B2(n25878), .C1(n16879), .C2(n25876), .A(
        n15002), .ZN(n14987) );
  OAI22_X2 U7144 ( .A1(n25873), .A2(n26537), .B1(n25871), .B2(n26633), .ZN(
        n15002) );
  NAND4_X2 U7145 ( .A1(n15005), .A2(n15006), .A3(n15007), .A4(n15008), .ZN(
        n14985) );
  AOI221_X2 U7146 ( .B1(n16860), .B2(n25870), .C1(n25867), .C2(n25422), .A(
        n15010), .ZN(n15008) );
  AOI221_X2 U7149 ( .B1(n25859), .B2(n25624), .C1(n25857), .C2(n25137), .A(
        n15016), .ZN(n15007) );
  OAI22_X2 U7150 ( .A1(n16891), .A2(n25856), .B1(n16863), .B2(n25853), .ZN(
        n15016) );
  AOI221_X2 U7153 ( .B1(n16883), .B2(n25852), .C1(n16874), .C2(n25850), .A(
        n15017), .ZN(n15006) );
  AOI221_X2 U7155 ( .B1(n16884), .B2(n25842), .C1(n16875), .C2(n25840), .A(
        n15018), .ZN(n15005) );
  OAI22_X2 U7156 ( .A1(n25838), .A2(n27145), .B1(n25835), .B2(n27209), .ZN(
        n15018) );
  NAND4_X2 U7159 ( .A1(n15024), .A2(n15025), .A3(n15026), .A4(n15027), .ZN(
        n15023) );
  AOI221_X2 U7160 ( .B1(n25906), .B2(n24973), .C1(n25903), .C2(n25421), .A(
        n15030), .ZN(n15027) );
  AOI221_X2 U7164 ( .B1(n25895), .B2(n24972), .C1(n25893), .C2(n25420), .A(
        n15035), .ZN(n15026) );
  OAI22_X2 U7165 ( .A1(n16849), .A2(n25891), .B1(n16821), .B2(n25889), .ZN(
        n15035) );
  AOI221_X2 U7168 ( .B1(n16834), .B2(n25888), .C1(n16825), .C2(n25886), .A(
        n15036), .ZN(n15025) );
  AOI221_X2 U7170 ( .B1(n16851), .B2(n25877), .C1(n16842), .C2(n25875), .A(
        n15039), .ZN(n15024) );
  OAI22_X2 U7171 ( .A1(n25874), .A2(n26538), .B1(n25871), .B2(n26634), .ZN(
        n15039) );
  NAND4_X2 U7172 ( .A1(n15042), .A2(n15043), .A3(n15044), .A4(n15045), .ZN(
        n15022) );
  AOI221_X2 U7173 ( .B1(n16823), .B2(n25869), .C1(n25868), .C2(n25419), .A(
        n15047), .ZN(n15045) );
  AOI221_X2 U7176 ( .B1(n25860), .B2(n25623), .C1(n25857), .C2(n25136), .A(
        n15053), .ZN(n15044) );
  OAI22_X2 U7177 ( .A1(n16854), .A2(n25855), .B1(n16826), .B2(n25853), .ZN(
        n15053) );
  AOI221_X2 U7180 ( .B1(n16846), .B2(n25851), .C1(n16837), .C2(n25849), .A(
        n15054), .ZN(n15043) );
  AOI221_X2 U7182 ( .B1(n16847), .B2(n25841), .C1(n16838), .C2(n25839), .A(
        n15055), .ZN(n15042) );
  OAI22_X2 U7183 ( .A1(n25837), .A2(n27146), .B1(n25836), .B2(n27210), .ZN(
        n15055) );
  NAND4_X2 U7186 ( .A1(n15061), .A2(n15062), .A3(n15063), .A4(n15064), .ZN(
        n15060) );
  AOI221_X2 U7187 ( .B1(n25905), .B2(n24971), .C1(n25904), .C2(n25418), .A(
        n15067), .ZN(n15064) );
  AOI221_X2 U7191 ( .B1(n25895), .B2(n24970), .C1(n25894), .C2(n25417), .A(
        n15072), .ZN(n15063) );
  OAI22_X2 U7192 ( .A1(n16812), .A2(n25892), .B1(n16784), .B2(n25889), .ZN(
        n15072) );
  AOI221_X2 U7195 ( .B1(n16797), .B2(n25887), .C1(n16788), .C2(n25885), .A(
        n15073), .ZN(n15062) );
  AOI221_X2 U7197 ( .B1(n16814), .B2(n25877), .C1(n16805), .C2(n25876), .A(
        n15076), .ZN(n15061) );
  OAI22_X2 U7198 ( .A1(n25873), .A2(n26539), .B1(n25871), .B2(n26635), .ZN(
        n15076) );
  NAND4_X2 U7199 ( .A1(n15079), .A2(n15080), .A3(n15081), .A4(n15082), .ZN(
        n15059) );
  AOI221_X2 U7200 ( .B1(n16786), .B2(n25870), .C1(n25868), .C2(n25416), .A(
        n15084), .ZN(n15082) );
  AOI221_X2 U7203 ( .B1(n25859), .B2(n25622), .C1(n25858), .C2(n25135), .A(
        n15090), .ZN(n15081) );
  OAI22_X2 U7204 ( .A1(n16817), .A2(n25855), .B1(n16789), .B2(n25853), .ZN(
        n15090) );
  AOI221_X2 U7207 ( .B1(n16809), .B2(n25851), .C1(n16800), .C2(n25850), .A(
        n15091), .ZN(n15080) );
  AOI221_X2 U7209 ( .B1(n16810), .B2(n25841), .C1(n16801), .C2(n25840), .A(
        n15092), .ZN(n15079) );
  OAI22_X2 U7210 ( .A1(n25838), .A2(n27147), .B1(n25835), .B2(n27211), .ZN(
        n15092) );
  NAND4_X2 U7213 ( .A1(n15098), .A2(n15099), .A3(n15100), .A4(n15101), .ZN(
        n15097) );
  AOI221_X2 U7214 ( .B1(n25906), .B2(n24969), .C1(n25904), .C2(n25415), .A(
        n15104), .ZN(n15101) );
  AOI221_X2 U7218 ( .B1(n25896), .B2(n24968), .C1(n25894), .C2(n25414), .A(
        n15109), .ZN(n15100) );
  OAI22_X2 U7219 ( .A1(n16775), .A2(n25891), .B1(n16747), .B2(n25890), .ZN(
        n15109) );
  AOI221_X2 U7222 ( .B1(n16760), .B2(n25887), .C1(n16751), .C2(n25886), .A(
        n15110), .ZN(n15099) );
  AOI221_X2 U7224 ( .B1(n16777), .B2(n25878), .C1(n16768), .C2(n25876), .A(
        n15113), .ZN(n15098) );
  OAI22_X2 U7225 ( .A1(n25873), .A2(n26540), .B1(n25872), .B2(n26636), .ZN(
        n15113) );
  NAND4_X2 U7226 ( .A1(n15116), .A2(n15117), .A3(n15118), .A4(n15119), .ZN(
        n15096) );
  AOI221_X2 U7227 ( .B1(n16749), .B2(n25869), .C1(n25868), .C2(n25413), .A(
        n15121), .ZN(n15119) );
  AOI221_X2 U7230 ( .B1(n25860), .B2(n24967), .C1(n25858), .C2(n25412), .A(
        n15127), .ZN(n15118) );
  OAI22_X2 U7231 ( .A1(n16780), .A2(n25856), .B1(n16752), .B2(n25854), .ZN(
        n15127) );
  AOI221_X2 U7234 ( .B1(n16772), .B2(n25852), .C1(n16763), .C2(n25850), .A(
        n15128), .ZN(n15117) );
  AOI221_X2 U7236 ( .B1(n16773), .B2(n25842), .C1(n16764), .C2(n25840), .A(
        n15129), .ZN(n15116) );
  OAI22_X2 U7237 ( .A1(n25838), .A2(n27148), .B1(n25836), .B2(n27212), .ZN(
        n15129) );
  OAI22_X2 U7238 ( .A1(n16744), .A2(n25907), .B1(n15132), .B2(n12153), .ZN(
        n23506) );
  NOR2_X2 U7239 ( .A1(n15133), .A2(n15134), .ZN(n15132) );
  NAND4_X2 U7240 ( .A1(n15135), .A2(n15136), .A3(n15137), .A4(n15138), .ZN(
        n15134) );
  AOI221_X2 U7241 ( .B1(n25906), .B2(n25621), .C1(n25904), .C2(n25134), .A(
        n15141), .ZN(n15138) );
  AOI221_X2 U7245 ( .B1(n25896), .B2(n25620), .C1(n25894), .C2(n25133), .A(
        n15146), .ZN(n15137) );
  OAI22_X2 U7246 ( .A1(n16738), .A2(n25891), .B1(n16710), .B2(n25890), .ZN(
        n15146) );
  AOI221_X2 U7249 ( .B1(n16723), .B2(n25888), .C1(n16714), .C2(n25886), .A(
        n15147), .ZN(n15136) );
  AOI221_X2 U7251 ( .B1(n16740), .B2(n25878), .C1(n16731), .C2(n25876), .A(
        n15150), .ZN(n15135) );
  OAI22_X2 U7252 ( .A1(n25873), .A2(n26541), .B1(n25872), .B2(n26637), .ZN(
        n15150) );
  NAND4_X2 U7253 ( .A1(n15153), .A2(n15154), .A3(n15155), .A4(n15156), .ZN(
        n15133) );
  AOI221_X2 U7254 ( .B1(n16712), .B2(n25869), .C1(n25868), .C2(n25411), .A(
        n15158), .ZN(n15156) );
  AOI221_X2 U7257 ( .B1(n25860), .B2(n25619), .C1(n25858), .C2(n25132), .A(
        n15164), .ZN(n15155) );
  OAI22_X2 U7258 ( .A1(n16743), .A2(n25855), .B1(n16715), .B2(n25854), .ZN(
        n15164) );
  AOI221_X2 U7261 ( .B1(n16735), .B2(n25852), .C1(n16726), .C2(n25850), .A(
        n15165), .ZN(n15154) );
  AOI221_X2 U7263 ( .B1(n16736), .B2(n25842), .C1(n16727), .C2(n25840), .A(
        n15166), .ZN(n15153) );
  OAI22_X2 U7264 ( .A1(n25838), .A2(n27149), .B1(n25836), .B2(n27213), .ZN(
        n15166) );
  OAI22_X2 U7265 ( .A1(n16707), .A2(n25907), .B1(n15169), .B2(n12153), .ZN(
        n23507) );
  NOR2_X2 U7266 ( .A1(n15170), .A2(n15171), .ZN(n15169) );
  NAND4_X2 U7267 ( .A1(n15172), .A2(n15173), .A3(n15174), .A4(n15175), .ZN(
        n15171) );
  AOI221_X2 U7268 ( .B1(n25906), .B2(n25618), .C1(n25904), .C2(n25131), .A(
        n15178), .ZN(n15175) );
  AOI221_X2 U7272 ( .B1(n25896), .B2(n25617), .C1(n25894), .C2(n25130), .A(
        n15183), .ZN(n15174) );
  OAI22_X2 U7273 ( .A1(n16701), .A2(n25891), .B1(n16673), .B2(n25889), .ZN(
        n15183) );
  AOI221_X2 U7276 ( .B1(n16686), .B2(n25888), .C1(n16677), .C2(n25886), .A(
        n15184), .ZN(n15173) );
  AOI221_X2 U7278 ( .B1(n16703), .B2(n25878), .C1(n16694), .C2(n25876), .A(
        n15187), .ZN(n15172) );
  OAI22_X2 U7279 ( .A1(n25873), .A2(n26542), .B1(n25872), .B2(n26638), .ZN(
        n15187) );
  NAND4_X2 U7280 ( .A1(n15190), .A2(n15191), .A3(n15192), .A4(n15193), .ZN(
        n15170) );
  AOI221_X2 U7281 ( .B1(n16675), .B2(n25869), .C1(n25868), .C2(n25410), .A(
        n15195), .ZN(n15193) );
  AOI221_X2 U7284 ( .B1(n25860), .B2(n25616), .C1(n25858), .C2(n25129), .A(
        n15201), .ZN(n15192) );
  OAI22_X2 U7285 ( .A1(n16706), .A2(n25855), .B1(n16678), .B2(n25853), .ZN(
        n15201) );
  AOI221_X2 U7288 ( .B1(n16698), .B2(n25852), .C1(n16689), .C2(n25850), .A(
        n15202), .ZN(n15191) );
  AOI221_X2 U7290 ( .B1(n16699), .B2(n25842), .C1(n16690), .C2(n25840), .A(
        n15203), .ZN(n15190) );
  OAI22_X2 U7291 ( .A1(n25838), .A2(n27150), .B1(n25836), .B2(n27214), .ZN(
        n15203) );
  OAI22_X2 U7292 ( .A1(n16670), .A2(n25907), .B1(n15206), .B2(n12153), .ZN(
        n23508) );
  NOR2_X2 U7293 ( .A1(n15207), .A2(n15208), .ZN(n15206) );
  NAND4_X2 U7294 ( .A1(n15209), .A2(n15210), .A3(n15211), .A4(n15212), .ZN(
        n15208) );
  AOI221_X2 U7295 ( .B1(n25906), .B2(n25615), .C1(n25904), .C2(n25128), .A(
        n15215), .ZN(n15212) );
  AOI221_X2 U7299 ( .B1(n25896), .B2(n25614), .C1(n25894), .C2(n25127), .A(
        n15220), .ZN(n15211) );
  OAI22_X2 U7300 ( .A1(n16664), .A2(n25892), .B1(n16636), .B2(n25890), .ZN(
        n15220) );
  AOI221_X2 U7303 ( .B1(n16649), .B2(n25888), .C1(n16640), .C2(n25886), .A(
        n15221), .ZN(n15210) );
  AOI221_X2 U7305 ( .B1(n16666), .B2(n25878), .C1(n16657), .C2(n25876), .A(
        n15224), .ZN(n15209) );
  OAI22_X2 U7306 ( .A1(n25874), .A2(n26543), .B1(n25871), .B2(n26639), .ZN(
        n15224) );
  NAND4_X2 U7307 ( .A1(n15227), .A2(n15228), .A3(n15229), .A4(n15230), .ZN(
        n15207) );
  AOI221_X2 U7308 ( .B1(n16638), .B2(n25869), .C1(n25868), .C2(n25409), .A(
        n15232), .ZN(n15230) );
  AOI221_X2 U7311 ( .B1(n25860), .B2(n25613), .C1(n25858), .C2(n25126), .A(
        n15238), .ZN(n15229) );
  OAI22_X2 U7312 ( .A1(n16669), .A2(n25856), .B1(n16641), .B2(n25853), .ZN(
        n15238) );
  AOI221_X2 U7315 ( .B1(n16661), .B2(n25852), .C1(n16652), .C2(n25850), .A(
        n15239), .ZN(n15228) );
  AOI221_X2 U7317 ( .B1(n16662), .B2(n25842), .C1(n16653), .C2(n25840), .A(
        n15240), .ZN(n15227) );
  OAI22_X2 U7318 ( .A1(n25837), .A2(n27151), .B1(n25836), .B2(n27215), .ZN(
        n15240) );
  OAI22_X2 U7319 ( .A1(n16633), .A2(n25909), .B1(n15243), .B2(n25908), .ZN(
        n23509) );
  NOR2_X2 U7320 ( .A1(n15244), .A2(n15245), .ZN(n15243) );
  NAND4_X2 U7321 ( .A1(n15246), .A2(n15247), .A3(n15248), .A4(n15249), .ZN(
        n15245) );
  AOI221_X2 U7322 ( .B1(n25906), .B2(n25612), .C1(n25904), .C2(n25125), .A(
        n15252), .ZN(n15249) );
  AOI221_X2 U7326 ( .B1(n25895), .B2(n25611), .C1(n25894), .C2(n25124), .A(
        n15257), .ZN(n15248) );
  OAI22_X2 U7327 ( .A1(n16627), .A2(n25892), .B1(n16599), .B2(n25890), .ZN(
        n15257) );
  AOI221_X2 U7330 ( .B1(n16612), .B2(n25888), .C1(n16603), .C2(n25885), .A(
        n15258), .ZN(n15247) );
  AOI221_X2 U7332 ( .B1(n16629), .B2(n25878), .C1(n16620), .C2(n25876), .A(
        n15261), .ZN(n15246) );
  OAI22_X2 U7333 ( .A1(n25874), .A2(n26544), .B1(n25871), .B2(n26640), .ZN(
        n15261) );
  NAND4_X2 U7334 ( .A1(n15264), .A2(n15265), .A3(n15266), .A4(n15267), .ZN(
        n15244) );
  AOI221_X2 U7335 ( .B1(n16601), .B2(n25869), .C1(n25868), .C2(n25408), .A(
        n15269), .ZN(n15267) );
  AOI221_X2 U7338 ( .B1(n25859), .B2(n25610), .C1(n25858), .C2(n25123), .A(
        n15275), .ZN(n15266) );
  OAI22_X2 U7339 ( .A1(n16632), .A2(n25856), .B1(n16604), .B2(n25853), .ZN(
        n15275) );
  AOI221_X2 U7342 ( .B1(n16624), .B2(n25852), .C1(n16615), .C2(n25850), .A(
        n15276), .ZN(n15265) );
  AOI221_X2 U7344 ( .B1(n16625), .B2(n25842), .C1(n16616), .C2(n25840), .A(
        n15277), .ZN(n15264) );
  OAI22_X2 U7345 ( .A1(n25837), .A2(n27152), .B1(n25835), .B2(n27216), .ZN(
        n15277) );
  OAI22_X2 U7346 ( .A1(n16596), .A2(n25907), .B1(n15280), .B2(n25908), .ZN(
        n23510) );
  NOR2_X2 U7347 ( .A1(n15281), .A2(n15282), .ZN(n15280) );
  NAND4_X2 U7348 ( .A1(n15283), .A2(n15284), .A3(n15285), .A4(n15286), .ZN(
        n15282) );
  AOI221_X2 U7349 ( .B1(n25905), .B2(n25609), .C1(n25904), .C2(n25122), .A(
        n15289), .ZN(n15286) );
  AOI221_X2 U7353 ( .B1(n25895), .B2(n25608), .C1(n25894), .C2(n25121), .A(
        n15294), .ZN(n15285) );
  OAI22_X2 U7354 ( .A1(n16590), .A2(n25891), .B1(n16562), .B2(n25889), .ZN(
        n15294) );
  AOI221_X2 U7357 ( .B1(n16575), .B2(n25888), .C1(n16566), .C2(n25885), .A(
        n15295), .ZN(n15284) );
  AOI221_X2 U7359 ( .B1(n16592), .B2(n25877), .C1(n16583), .C2(n25876), .A(
        n15298), .ZN(n15283) );
  OAI22_X2 U7360 ( .A1(n25873), .A2(n26545), .B1(n25871), .B2(n26641), .ZN(
        n15298) );
  NAND4_X2 U7361 ( .A1(n15301), .A2(n15302), .A3(n15303), .A4(n15304), .ZN(
        n15281) );
  AOI221_X2 U7362 ( .B1(n16564), .B2(n25870), .C1(n25868), .C2(n25407), .A(
        n15306), .ZN(n15304) );
  AOI221_X2 U7365 ( .B1(n25859), .B2(n25607), .C1(n25858), .C2(n25120), .A(
        n15312), .ZN(n15303) );
  OAI22_X2 U7366 ( .A1(n16595), .A2(n25855), .B1(n16567), .B2(n25854), .ZN(
        n15312) );
  AOI221_X2 U7369 ( .B1(n16587), .B2(n25851), .C1(n16578), .C2(n25850), .A(
        n15313), .ZN(n15302) );
  AOI221_X2 U7371 ( .B1(n16588), .B2(n25841), .C1(n16579), .C2(n25840), .A(
        n15314), .ZN(n15301) );
  OAI22_X2 U7372 ( .A1(n25838), .A2(n27153), .B1(n25835), .B2(n27217), .ZN(
        n15314) );
  OAI22_X2 U7373 ( .A1(n16559), .A2(n25907), .B1(n15317), .B2(n12153), .ZN(
        n23511) );
  NOR2_X2 U7374 ( .A1(n15318), .A2(n15319), .ZN(n15317) );
  NAND4_X2 U7375 ( .A1(n15320), .A2(n15321), .A3(n15322), .A4(n15323), .ZN(
        n15319) );
  AOI221_X2 U7376 ( .B1(n25906), .B2(n25606), .C1(n25904), .C2(n25119), .A(
        n15326), .ZN(n15323) );
  AOI221_X2 U7380 ( .B1(n25896), .B2(n25605), .C1(n25894), .C2(n25118), .A(
        n15331), .ZN(n15322) );
  OAI22_X2 U7381 ( .A1(n16553), .A2(n25892), .B1(n16525), .B2(n25889), .ZN(
        n15331) );
  AOI221_X2 U7384 ( .B1(n16538), .B2(n25888), .C1(n16529), .C2(n25886), .A(
        n15332), .ZN(n15321) );
  AOI221_X2 U7386 ( .B1(n16555), .B2(n25878), .C1(n16546), .C2(n25876), .A(
        n15335), .ZN(n15320) );
  OAI22_X2 U7387 ( .A1(n25874), .A2(n26546), .B1(n25871), .B2(n26642), .ZN(
        n15335) );
  NAND4_X2 U7388 ( .A1(n15338), .A2(n15339), .A3(n15340), .A4(n15341), .ZN(
        n15318) );
  AOI221_X2 U7389 ( .B1(n16527), .B2(n25869), .C1(n25868), .C2(n25406), .A(
        n15343), .ZN(n15341) );
  AOI221_X2 U7392 ( .B1(n25860), .B2(n25604), .C1(n25858), .C2(n25117), .A(
        n15349), .ZN(n15340) );
  OAI22_X2 U7393 ( .A1(n16558), .A2(n25856), .B1(n16530), .B2(n25854), .ZN(
        n15349) );
  AOI221_X2 U7396 ( .B1(n16550), .B2(n25852), .C1(n16541), .C2(n25850), .A(
        n15350), .ZN(n15339) );
  AOI221_X2 U7398 ( .B1(n16551), .B2(n25842), .C1(n16542), .C2(n25840), .A(
        n15351), .ZN(n15338) );
  OAI22_X2 U7399 ( .A1(n25837), .A2(n27154), .B1(n25836), .B2(n27218), .ZN(
        n15351) );
  OAI22_X2 U7400 ( .A1(n16522), .A2(n25907), .B1(n15354), .B2(n12153), .ZN(
        n23512) );
  NOR2_X2 U7401 ( .A1(n15355), .A2(n15356), .ZN(n15354) );
  NAND4_X2 U7402 ( .A1(n15357), .A2(n15358), .A3(n15359), .A4(n15360), .ZN(
        n15356) );
  AOI221_X2 U7403 ( .B1(n25906), .B2(n25603), .C1(n25904), .C2(n25116), .A(
        n15363), .ZN(n15360) );
  AOI221_X2 U7407 ( .B1(n25895), .B2(n25602), .C1(n25894), .C2(n25115), .A(
        n15368), .ZN(n15359) );
  OAI22_X2 U7408 ( .A1(n16516), .A2(n25892), .B1(n16488), .B2(n25890), .ZN(
        n15368) );
  AOI221_X2 U7411 ( .B1(n16501), .B2(n25888), .C1(n16492), .C2(n25885), .A(
        n15369), .ZN(n15358) );
  AOI221_X2 U7413 ( .B1(n16518), .B2(n25878), .C1(n16509), .C2(n25876), .A(
        n15372), .ZN(n15357) );
  OAI22_X2 U7414 ( .A1(n25874), .A2(n26547), .B1(n25872), .B2(n26643), .ZN(
        n15372) );
  NAND4_X2 U7415 ( .A1(n15375), .A2(n15376), .A3(n15377), .A4(n15378), .ZN(
        n15355) );
  AOI221_X2 U7416 ( .B1(n16490), .B2(n25869), .C1(n25868), .C2(n25405), .A(
        n15380), .ZN(n15378) );
  AOI221_X2 U7419 ( .B1(n25859), .B2(n25601), .C1(n25858), .C2(n25114), .A(
        n15386), .ZN(n15377) );
  OAI22_X2 U7420 ( .A1(n16521), .A2(n25856), .B1(n16493), .B2(n25854), .ZN(
        n15386) );
  AOI221_X2 U7423 ( .B1(n16513), .B2(n25852), .C1(n16504), .C2(n25850), .A(
        n15387), .ZN(n15376) );
  AOI221_X2 U7425 ( .B1(n16514), .B2(n25842), .C1(n16505), .C2(n25840), .A(
        n15388), .ZN(n15375) );
  OAI22_X2 U7426 ( .A1(n25838), .A2(n27155), .B1(n25836), .B2(n27219), .ZN(
        n15388) );
  OAI22_X2 U7427 ( .A1(n16485), .A2(n25907), .B1(n15391), .B2(n12153), .ZN(
        n23513) );
  NOR2_X2 U7428 ( .A1(n15392), .A2(n15393), .ZN(n15391) );
  NAND4_X2 U7429 ( .A1(n15394), .A2(n15395), .A3(n15396), .A4(n15397), .ZN(
        n15393) );
  AOI221_X2 U7430 ( .B1(n25905), .B2(n25600), .C1(n25904), .C2(n25113), .A(
        n15400), .ZN(n15397) );
  AOI221_X2 U7434 ( .B1(n25895), .B2(n25599), .C1(n25894), .C2(n25112), .A(
        n15405), .ZN(n15396) );
  OAI22_X2 U7435 ( .A1(n16479), .A2(n25892), .B1(n16451), .B2(n25890), .ZN(
        n15405) );
  AOI221_X2 U7438 ( .B1(n16464), .B2(n25887), .C1(n16455), .C2(n25885), .A(
        n15406), .ZN(n15395) );
  AOI221_X2 U7440 ( .B1(n16481), .B2(n25877), .C1(n16472), .C2(n25876), .A(
        n15409), .ZN(n15394) );
  OAI22_X2 U7441 ( .A1(n25874), .A2(n26548), .B1(n25872), .B2(n26644), .ZN(
        n15409) );
  NAND4_X2 U7442 ( .A1(n15412), .A2(n15413), .A3(n15414), .A4(n15415), .ZN(
        n15392) );
  AOI221_X2 U7443 ( .B1(n16453), .B2(n25870), .C1(n25868), .C2(n25404), .A(
        n15417), .ZN(n15415) );
  AOI221_X2 U7446 ( .B1(n25859), .B2(n25598), .C1(n25858), .C2(n25111), .A(
        n15423), .ZN(n15414) );
  OAI22_X2 U7447 ( .A1(n16484), .A2(n25856), .B1(n16456), .B2(n25854), .ZN(
        n15423) );
  AOI221_X2 U7450 ( .B1(n16476), .B2(n25851), .C1(n16467), .C2(n25850), .A(
        n15424), .ZN(n15413) );
  AOI221_X2 U7452 ( .B1(n16477), .B2(n25841), .C1(n16468), .C2(n25840), .A(
        n15425), .ZN(n15412) );
  OAI22_X2 U7453 ( .A1(n25837), .A2(n27156), .B1(n25836), .B2(n27220), .ZN(
        n15425) );
  OAI22_X2 U7454 ( .A1(n16448), .A2(n25909), .B1(n15428), .B2(n12153), .ZN(
        n23514) );
  NOR2_X2 U7455 ( .A1(n15429), .A2(n15430), .ZN(n15428) );
  NAND4_X2 U7456 ( .A1(n15431), .A2(n15432), .A3(n15433), .A4(n15434), .ZN(
        n15430) );
  AOI221_X2 U7457 ( .B1(n25905), .B2(n25597), .C1(n25904), .C2(n25110), .A(
        n15437), .ZN(n15434) );
  AOI221_X2 U7461 ( .B1(n25895), .B2(n25596), .C1(n25894), .C2(n25109), .A(
        n15442), .ZN(n15433) );
  OAI22_X2 U7462 ( .A1(n16442), .A2(n25892), .B1(n16414), .B2(n25890), .ZN(
        n15442) );
  AOI221_X2 U7465 ( .B1(n16427), .B2(n25888), .C1(n16418), .C2(n25886), .A(
        n15443), .ZN(n15432) );
  AOI221_X2 U7467 ( .B1(n16444), .B2(n25877), .C1(n16435), .C2(n25876), .A(
        n15446), .ZN(n15431) );
  OAI22_X2 U7468 ( .A1(n25873), .A2(n26549), .B1(n25872), .B2(n26645), .ZN(
        n15446) );
  NAND4_X2 U7469 ( .A1(n15449), .A2(n15450), .A3(n15451), .A4(n15452), .ZN(
        n15429) );
  AOI221_X2 U7470 ( .B1(n16416), .B2(n25870), .C1(n25868), .C2(n25403), .A(
        n15454), .ZN(n15452) );
  AOI221_X2 U7473 ( .B1(n25859), .B2(n25595), .C1(n25858), .C2(n25108), .A(
        n15460), .ZN(n15451) );
  OAI22_X2 U7474 ( .A1(n16447), .A2(n25856), .B1(n16419), .B2(n25854), .ZN(
        n15460) );
  AOI221_X2 U7477 ( .B1(n16439), .B2(n25851), .C1(n16430), .C2(n25850), .A(
        n15461), .ZN(n15450) );
  AOI221_X2 U7479 ( .B1(n16440), .B2(n25841), .C1(n16431), .C2(n25840), .A(
        n15462), .ZN(n15449) );
  OAI22_X2 U7480 ( .A1(n25838), .A2(n27157), .B1(n25836), .B2(n27221), .ZN(
        n15462) );
  OAI22_X2 U7481 ( .A1(n16411), .A2(n25909), .B1(n15465), .B2(n12153), .ZN(
        n23515) );
  NOR2_X2 U7482 ( .A1(n15466), .A2(n15467), .ZN(n15465) );
  NAND4_X2 U7483 ( .A1(n15468), .A2(n15469), .A3(n15470), .A4(n15471), .ZN(
        n15467) );
  AOI221_X2 U7484 ( .B1(n25905), .B2(n25594), .C1(n25904), .C2(n25107), .A(
        n15474), .ZN(n15471) );
  AOI221_X2 U7493 ( .B1(n25896), .B2(n25593), .C1(n25894), .C2(n25106), .A(
        n15483), .ZN(n15470) );
  OAI22_X2 U7494 ( .A1(n16405), .A2(n25891), .B1(n16377), .B2(n25890), .ZN(
        n15483) );
  AOI221_X2 U7502 ( .B1(n16390), .B2(n25888), .C1(n16381), .C2(n25885), .A(
        n15485), .ZN(n15469) );
  AOI221_X2 U7510 ( .B1(n16407), .B2(n25877), .C1(n16398), .C2(n25876), .A(
        n15489), .ZN(n15468) );
  OAI22_X2 U7511 ( .A1(n25873), .A2(n26550), .B1(n25872), .B2(n26646), .ZN(
        n15489) );
  NAND4_X2 U7516 ( .A1(n15492), .A2(n15493), .A3(n15494), .A4(n15495), .ZN(
        n15466) );
  AOI221_X2 U7517 ( .B1(n16379), .B2(n25870), .C1(n25868), .C2(n25402), .A(
        n15497), .ZN(n15495) );
  AOI221_X2 U7525 ( .B1(n25860), .B2(n25592), .C1(n25858), .C2(n25105), .A(
        n15503), .ZN(n15494) );
  OAI22_X2 U7526 ( .A1(n16410), .A2(n25855), .B1(n16382), .B2(n25854), .ZN(
        n15503) );
  AOI221_X2 U7533 ( .B1(n16402), .B2(n25851), .C1(n16393), .C2(n25850), .A(
        n15504), .ZN(n15493) );
  AOI221_X2 U7540 ( .B1(n16403), .B2(n25841), .C1(n16394), .C2(n25840), .A(
        n15505), .ZN(n15492) );
  OAI22_X2 U7541 ( .A1(n25837), .A2(n27158), .B1(n25836), .B2(n27222), .ZN(
        n15505) );
  NAND2_X2 U7544 ( .A1(n27803), .A2(n15509), .ZN(n12840) );
  NAND2_X2 U7545 ( .A1(n27802), .A2(n15509), .ZN(n12831) );
  NAND2_X2 U7546 ( .A1(n15511), .A2(n15509), .ZN(n12827) );
  NAND2_X2 U7549 ( .A1(n27803), .A2(n27804), .ZN(n12841) );
  NAND2_X2 U7550 ( .A1(n27802), .A2(n27804), .ZN(n12832) );
  NAND2_X2 U7551 ( .A1(n15511), .A2(n27804), .ZN(n12828) );
  NAND2_X2 U7552 ( .A1(n27804), .A2(n15513), .ZN(n12816) );
  NAND2_X2 U7556 ( .A1(n27803), .A2(n15515), .ZN(n12839) );
  NAND2_X2 U7557 ( .A1(n27802), .A2(n15515), .ZN(n12830) );
  NAND2_X2 U7558 ( .A1(n15511), .A2(n15515), .ZN(n12826) );
  NAND2_X2 U7559 ( .A1(n15515), .A2(n15513), .ZN(n12815) );
  NAND2_X2 U7563 ( .A1(n27803), .A2(n15516), .ZN(n12838) );
  NAND2_X2 U7565 ( .A1(n27802), .A2(n15516), .ZN(n12829) );
  NAND2_X2 U7567 ( .A1(n15511), .A2(n15516), .ZN(n12825) );
  NOR2_X2 U7568 ( .A1(n25245), .A2(n24890), .ZN(n15511) );
  NAND2_X2 U7569 ( .A1(n15516), .A2(n15513), .ZN(n12814) );
  NOR2_X2 U7570 ( .A1(n22395), .A2(n22396), .ZN(n15516) );
  NAND4_X2 U7573 ( .A1(n15484), .A2(n15488), .A3(n15522), .A4(n15523), .ZN(
        n15521) );
  NOR4_X2 U7574 ( .A1(n12799), .A2(n12803), .A3(n12811), .A4(n12788), .ZN(
        n15523) );
  NOR3_X2 U7578 ( .A1(add_180_A_1_), .A2(n22394), .A3(add_180_A_3_), .ZN(
        n15526) );
  NOR3_X2 U7580 ( .A1(n12812), .A2(n12813), .A3(n12786), .ZN(n15522) );
  NAND3_X2 U7583 ( .A1(n22392), .A2(n22394), .A3(n25250), .ZN(n15484) );
  NAND2_X2 U7585 ( .A1(n15513), .A2(n15509), .ZN(n12817) );
  NOR2_X2 U7586 ( .A1(n25246), .A2(n22396), .ZN(n15509) );
  NAND2_X2 U7587 ( .A1(n22396), .A2(n25246), .ZN(n15514) );
  OAI22_X2 U7589 ( .A1(n22396), .A2(n26286), .B1(n15531), .B2(n15534), .ZN(
        n23517) );
  NOR2_X2 U7593 ( .A1(n22398), .A2(n22397), .ZN(n15513) );
  NAND2_X2 U7595 ( .A1(n22398), .A2(n25245), .ZN(n15517) );
  NAND2_X2 U7597 ( .A1(n22397), .A2(n24890), .ZN(n15518) );
  OAI22_X2 U7598 ( .A1(n22398), .A2(n15536), .B1(n24890), .B2(n15531), .ZN(
        n23519) );
  NAND2_X2 U7600 ( .A1(n12813), .A2(n11634), .ZN(n15530) );
  NOR2_X2 U7602 ( .A1(n15537), .A2(n15538), .ZN(n15536) );
  OAI22_X2 U7603 ( .A1(n15488), .A2(n15539), .B1(n22391), .B2(n15540), .ZN(
        n23520) );
  NAND3_X2 U7605 ( .A1(add_180_A_0_), .A2(add_180_A_2_), .A3(n25250), .ZN(
        n15488) );
  OAI22_X2 U7613 ( .A1(n22393), .A2(n15545), .B1(n15539), .B2(n15546), .ZN(
        n23522) );
  OAI22_X2 U7616 ( .A1(n22394), .A2(n26287), .B1(add_180_A_0_), .B2(n15539), 
        .ZN(n23523) );
  NAND2_X2 U7617 ( .A1(n15538), .A2(n26287), .ZN(n15539) );
  NOR2_X2 U7618 ( .A1(n26293), .A2(n12813), .ZN(n15538) );
  NOR2_X2 U7624 ( .A1(n26293), .A2(n13093), .ZN(n15537) );
  NOR2_X2 U7625 ( .A1(n16374), .A2(n22381), .ZN(n13093) );
  OAI22_X2 U7626 ( .A1(n26382), .A2(n26551), .B1(n25833), .B2(n15550), .ZN(
        n23524) );
  OAI22_X2 U7628 ( .A1(n26382), .A2(n26552), .B1(n25827), .B2(n15550), .ZN(
        n23525) );
  OAI22_X2 U7630 ( .A1(n26382), .A2(n26553), .B1(n25825), .B2(n15550), .ZN(
        n23526) );
  OAI22_X2 U7632 ( .A1(n26382), .A2(n26554), .B1(n25822), .B2(n15550), .ZN(
        n23527) );
  OAI22_X2 U7634 ( .A1(n26382), .A2(n26555), .B1(n25819), .B2(n15550), .ZN(
        n23528) );
  OAI22_X2 U7636 ( .A1(n26382), .A2(n26556), .B1(n25816), .B2(n15550), .ZN(
        n23529) );
  OAI22_X2 U7638 ( .A1(n26382), .A2(n26557), .B1(n25813), .B2(n15550), .ZN(
        n23530) );
  OAI22_X2 U7640 ( .A1(n26382), .A2(n26558), .B1(n25810), .B2(n15550), .ZN(
        n23531) );
  OAI22_X2 U7642 ( .A1(n26382), .A2(n26559), .B1(n25807), .B2(n15550), .ZN(
        n23532) );
  OAI22_X2 U7644 ( .A1(n26382), .A2(n26560), .B1(n25804), .B2(n15550), .ZN(
        n23533) );
  OAI22_X2 U7646 ( .A1(n26382), .A2(n26561), .B1(n25801), .B2(n15550), .ZN(
        n23534) );
  OAI22_X2 U7648 ( .A1(n26382), .A2(n26562), .B1(n25796), .B2(n15550), .ZN(
        n23535) );
  OAI22_X2 U7650 ( .A1(n26382), .A2(n26563), .B1(n25791), .B2(n15550), .ZN(
        n23536) );
  OAI22_X2 U7652 ( .A1(n26382), .A2(n26564), .B1(n25789), .B2(n15550), .ZN(
        n23537) );
  OAI22_X2 U7654 ( .A1(n26382), .A2(n26565), .B1(n25786), .B2(n15550), .ZN(
        n23538) );
  OAI22_X2 U7656 ( .A1(n26382), .A2(n26566), .B1(n25783), .B2(n15550), .ZN(
        n23539) );
  OAI22_X2 U7660 ( .A1(n26381), .A2(n27543), .B1(n25833), .B2(n15567), .ZN(
        n23540) );
  OAI22_X2 U7662 ( .A1(n26381), .A2(n27544), .B1(n25828), .B2(n15567), .ZN(
        n23541) );
  OAI22_X2 U7664 ( .A1(n26381), .A2(n27545), .B1(n25825), .B2(n15567), .ZN(
        n23542) );
  OAI22_X2 U7666 ( .A1(n26381), .A2(n27546), .B1(n25822), .B2(n15567), .ZN(
        n23543) );
  OAI22_X2 U7668 ( .A1(n26381), .A2(n27547), .B1(n25819), .B2(n15567), .ZN(
        n23544) );
  OAI22_X2 U7670 ( .A1(n26381), .A2(n27548), .B1(n25816), .B2(n15567), .ZN(
        n23545) );
  OAI22_X2 U7672 ( .A1(n26381), .A2(n27549), .B1(n25813), .B2(n15567), .ZN(
        n23546) );
  OAI22_X2 U7674 ( .A1(n26381), .A2(n27550), .B1(n25810), .B2(n15567), .ZN(
        n23547) );
  OAI22_X2 U7676 ( .A1(n26381), .A2(n27551), .B1(n25807), .B2(n15567), .ZN(
        n23548) );
  OAI22_X2 U7678 ( .A1(n26381), .A2(n27552), .B1(n25804), .B2(n15567), .ZN(
        n23549) );
  OAI22_X2 U7680 ( .A1(n26381), .A2(n27553), .B1(n25801), .B2(n15567), .ZN(
        n23550) );
  OAI22_X2 U7682 ( .A1(n26381), .A2(n27554), .B1(n25797), .B2(n15567), .ZN(
        n23551) );
  OAI22_X2 U7684 ( .A1(n26381), .A2(n27555), .B1(n25792), .B2(n15567), .ZN(
        n23552) );
  OAI22_X2 U7686 ( .A1(n26381), .A2(n27556), .B1(n25789), .B2(n15567), .ZN(
        n23553) );
  OAI22_X2 U7688 ( .A1(n26381), .A2(n27557), .B1(n25786), .B2(n15567), .ZN(
        n23554) );
  OAI22_X2 U7690 ( .A1(n26381), .A2(n27558), .B1(n25783), .B2(n15567), .ZN(
        n23555) );
  OAI22_X2 U7694 ( .A1(n26380), .A2(n26775), .B1(n25834), .B2(n15569), .ZN(
        n23556) );
  OAI22_X2 U7696 ( .A1(n26380), .A2(n26776), .B1(n25828), .B2(n15569), .ZN(
        n23557) );
  OAI22_X2 U7698 ( .A1(n26380), .A2(n26777), .B1(n25826), .B2(n15569), .ZN(
        n23558) );
  OAI22_X2 U7700 ( .A1(n26380), .A2(n26778), .B1(n25823), .B2(n15569), .ZN(
        n23559) );
  OAI22_X2 U7702 ( .A1(n26380), .A2(n26779), .B1(n25820), .B2(n15569), .ZN(
        n23560) );
  OAI22_X2 U7704 ( .A1(n26380), .A2(n26780), .B1(n25817), .B2(n15569), .ZN(
        n23561) );
  OAI22_X2 U7706 ( .A1(n26380), .A2(n26781), .B1(n25814), .B2(n15569), .ZN(
        n23562) );
  OAI22_X2 U7708 ( .A1(n26380), .A2(n26782), .B1(n25811), .B2(n15569), .ZN(
        n23563) );
  OAI22_X2 U7710 ( .A1(n26380), .A2(n26783), .B1(n25808), .B2(n15569), .ZN(
        n23564) );
  OAI22_X2 U7712 ( .A1(n26380), .A2(n26784), .B1(n25805), .B2(n15569), .ZN(
        n23565) );
  OAI22_X2 U7714 ( .A1(n26380), .A2(n26785), .B1(n25802), .B2(n15569), .ZN(
        n23566) );
  OAI22_X2 U7716 ( .A1(n26380), .A2(n26786), .B1(n25797), .B2(n15569), .ZN(
        n23567) );
  OAI22_X2 U7718 ( .A1(n26380), .A2(n26787), .B1(n25792), .B2(n15569), .ZN(
        n23568) );
  OAI22_X2 U7720 ( .A1(n26380), .A2(n26788), .B1(n25790), .B2(n15569), .ZN(
        n23569) );
  OAI22_X2 U7722 ( .A1(n26380), .A2(n26789), .B1(n25787), .B2(n15569), .ZN(
        n23570) );
  OAI22_X2 U7724 ( .A1(n26380), .A2(n26790), .B1(n25784), .B2(n15569), .ZN(
        n23571) );
  OAI22_X2 U7728 ( .A1(n26379), .A2(n27031), .B1(n25832), .B2(n15572), .ZN(
        n23572) );
  OAI22_X2 U7730 ( .A1(n26379), .A2(n27032), .B1(n25828), .B2(n15572), .ZN(
        n23573) );
  OAI22_X2 U7732 ( .A1(n26379), .A2(n27033), .B1(n25824), .B2(n15572), .ZN(
        n23574) );
  OAI22_X2 U7734 ( .A1(n26379), .A2(n27034), .B1(n25821), .B2(n15572), .ZN(
        n23575) );
  OAI22_X2 U7736 ( .A1(n26379), .A2(n27035), .B1(n25818), .B2(n15572), .ZN(
        n23576) );
  OAI22_X2 U7738 ( .A1(n26379), .A2(n27036), .B1(n25815), .B2(n15572), .ZN(
        n23577) );
  OAI22_X2 U7740 ( .A1(n26379), .A2(n27037), .B1(n25812), .B2(n15572), .ZN(
        n23578) );
  OAI22_X2 U7742 ( .A1(n26379), .A2(n27038), .B1(n25809), .B2(n15572), .ZN(
        n23579) );
  OAI22_X2 U7744 ( .A1(n26379), .A2(n27039), .B1(n25806), .B2(n15572), .ZN(
        n23580) );
  OAI22_X2 U7746 ( .A1(n26379), .A2(n27040), .B1(n25803), .B2(n15572), .ZN(
        n23581) );
  OAI22_X2 U7748 ( .A1(n26379), .A2(n27041), .B1(n25800), .B2(n15572), .ZN(
        n23582) );
  OAI22_X2 U7750 ( .A1(n26379), .A2(n27042), .B1(n25797), .B2(n15572), .ZN(
        n23583) );
  OAI22_X2 U7752 ( .A1(n26379), .A2(n27043), .B1(n25792), .B2(n15572), .ZN(
        n23584) );
  OAI22_X2 U7754 ( .A1(n26379), .A2(n27044), .B1(n25788), .B2(n15572), .ZN(
        n23585) );
  OAI22_X2 U7756 ( .A1(n26379), .A2(n27045), .B1(n25785), .B2(n15572), .ZN(
        n23586) );
  OAI22_X2 U7758 ( .A1(n26379), .A2(n27046), .B1(n25782), .B2(n15572), .ZN(
        n23587) );
  OAI22_X2 U7762 ( .A1(n26378), .A2(n27287), .B1(n25832), .B2(n15590), .ZN(
        n23588) );
  OAI22_X2 U7764 ( .A1(n26378), .A2(n27288), .B1(n25828), .B2(n15590), .ZN(
        n23589) );
  OAI22_X2 U7766 ( .A1(n26378), .A2(n27289), .B1(n25824), .B2(n15590), .ZN(
        n23590) );
  OAI22_X2 U7768 ( .A1(n26378), .A2(n27290), .B1(n25821), .B2(n15590), .ZN(
        n23591) );
  OAI22_X2 U7770 ( .A1(n26378), .A2(n27291), .B1(n25818), .B2(n15590), .ZN(
        n23592) );
  OAI22_X2 U7772 ( .A1(n26378), .A2(n27292), .B1(n25815), .B2(n15590), .ZN(
        n23593) );
  OAI22_X2 U7774 ( .A1(n26378), .A2(n27293), .B1(n25812), .B2(n15590), .ZN(
        n23594) );
  OAI22_X2 U7776 ( .A1(n26378), .A2(n27294), .B1(n25809), .B2(n15590), .ZN(
        n23595) );
  OAI22_X2 U7778 ( .A1(n26378), .A2(n27295), .B1(n25806), .B2(n15590), .ZN(
        n23596) );
  OAI22_X2 U7780 ( .A1(n26378), .A2(n27296), .B1(n25803), .B2(n15590), .ZN(
        n23597) );
  OAI22_X2 U7782 ( .A1(n26378), .A2(n27297), .B1(n25800), .B2(n15590), .ZN(
        n23598) );
  OAI22_X2 U7784 ( .A1(n26378), .A2(n27298), .B1(n25797), .B2(n15590), .ZN(
        n23599) );
  OAI22_X2 U7786 ( .A1(n26378), .A2(n27299), .B1(n25792), .B2(n15590), .ZN(
        n23600) );
  OAI22_X2 U7788 ( .A1(n26378), .A2(n27300), .B1(n25788), .B2(n15590), .ZN(
        n23601) );
  OAI22_X2 U7790 ( .A1(n26378), .A2(n27301), .B1(n25785), .B2(n15590), .ZN(
        n23602) );
  OAI22_X2 U7792 ( .A1(n26378), .A2(n27302), .B1(n25782), .B2(n15590), .ZN(
        n23603) );
  OAI22_X2 U7797 ( .A1(n26373), .A2(n26711), .B1(n25833), .B2(n15609), .ZN(
        n23604) );
  OAI22_X2 U7799 ( .A1(n26373), .A2(n26712), .B1(n25828), .B2(n15609), .ZN(
        n23605) );
  OAI22_X2 U7801 ( .A1(n26373), .A2(n26713), .B1(n25825), .B2(n15609), .ZN(
        n23606) );
  OAI22_X2 U7803 ( .A1(n26373), .A2(n26714), .B1(n25822), .B2(n15609), .ZN(
        n23607) );
  OAI22_X2 U7805 ( .A1(n26373), .A2(n26715), .B1(n25819), .B2(n15609), .ZN(
        n23608) );
  OAI22_X2 U7807 ( .A1(n26373), .A2(n26716), .B1(n25816), .B2(n15609), .ZN(
        n23609) );
  OAI22_X2 U7809 ( .A1(n26373), .A2(n26717), .B1(n25813), .B2(n15609), .ZN(
        n23610) );
  OAI22_X2 U7811 ( .A1(n26373), .A2(n26718), .B1(n25810), .B2(n15609), .ZN(
        n23611) );
  OAI22_X2 U7813 ( .A1(n26373), .A2(n26719), .B1(n25807), .B2(n15609), .ZN(
        n23612) );
  OAI22_X2 U7815 ( .A1(n26373), .A2(n26720), .B1(n25804), .B2(n15609), .ZN(
        n23613) );
  OAI22_X2 U7817 ( .A1(n26373), .A2(n26721), .B1(n25801), .B2(n15609), .ZN(
        n23614) );
  OAI22_X2 U7819 ( .A1(n26373), .A2(n26722), .B1(n25797), .B2(n15609), .ZN(
        n23615) );
  OAI22_X2 U7821 ( .A1(n26373), .A2(n26723), .B1(n25792), .B2(n15609), .ZN(
        n23616) );
  OAI22_X2 U7823 ( .A1(n26373), .A2(n26724), .B1(n25789), .B2(n15609), .ZN(
        n23617) );
  OAI22_X2 U7825 ( .A1(n26373), .A2(n26725), .B1(n25786), .B2(n15609), .ZN(
        n23618) );
  OAI22_X2 U7827 ( .A1(n26373), .A2(n26726), .B1(n25783), .B2(n15609), .ZN(
        n23619) );
  OAI22_X2 U7831 ( .A1(n26372), .A2(n27559), .B1(n25834), .B2(n15626), .ZN(
        n23620) );
  OAI22_X2 U7833 ( .A1(n26372), .A2(n27560), .B1(n25828), .B2(n15626), .ZN(
        n23621) );
  OAI22_X2 U7835 ( .A1(n26372), .A2(n27561), .B1(n25826), .B2(n15626), .ZN(
        n23622) );
  OAI22_X2 U7837 ( .A1(n26372), .A2(n27562), .B1(n25823), .B2(n15626), .ZN(
        n23623) );
  OAI22_X2 U7839 ( .A1(n26372), .A2(n27563), .B1(n25820), .B2(n15626), .ZN(
        n23624) );
  OAI22_X2 U7841 ( .A1(n26372), .A2(n27564), .B1(n25817), .B2(n15626), .ZN(
        n23625) );
  OAI22_X2 U7843 ( .A1(n26372), .A2(n27565), .B1(n25814), .B2(n15626), .ZN(
        n23626) );
  OAI22_X2 U7845 ( .A1(n26372), .A2(n27566), .B1(n25811), .B2(n15626), .ZN(
        n23627) );
  OAI22_X2 U7847 ( .A1(n26372), .A2(n27567), .B1(n25808), .B2(n15626), .ZN(
        n23628) );
  OAI22_X2 U7849 ( .A1(n26372), .A2(n27568), .B1(n25805), .B2(n15626), .ZN(
        n23629) );
  OAI22_X2 U7851 ( .A1(n26372), .A2(n27569), .B1(n25802), .B2(n15626), .ZN(
        n23630) );
  OAI22_X2 U7853 ( .A1(n26372), .A2(n27570), .B1(n25797), .B2(n15626), .ZN(
        n23631) );
  OAI22_X2 U7855 ( .A1(n26372), .A2(n27571), .B1(n25792), .B2(n15626), .ZN(
        n23632) );
  OAI22_X2 U7857 ( .A1(n26372), .A2(n27572), .B1(n25790), .B2(n15626), .ZN(
        n23633) );
  OAI22_X2 U7859 ( .A1(n26372), .A2(n27573), .B1(n25787), .B2(n15626), .ZN(
        n23634) );
  OAI22_X2 U7861 ( .A1(n26372), .A2(n27574), .B1(n25784), .B2(n15626), .ZN(
        n23635) );
  OAI22_X2 U7865 ( .A1(n26371), .A2(n26791), .B1(n25834), .B2(n15628), .ZN(
        n23636) );
  OAI22_X2 U7867 ( .A1(n26371), .A2(n26792), .B1(n25828), .B2(n15628), .ZN(
        n23637) );
  OAI22_X2 U7869 ( .A1(n26371), .A2(n26793), .B1(n25826), .B2(n15628), .ZN(
        n23638) );
  OAI22_X2 U7871 ( .A1(n26371), .A2(n26794), .B1(n25823), .B2(n15628), .ZN(
        n23639) );
  OAI22_X2 U7873 ( .A1(n26371), .A2(n26795), .B1(n25820), .B2(n15628), .ZN(
        n23640) );
  OAI22_X2 U7875 ( .A1(n26371), .A2(n26796), .B1(n25817), .B2(n15628), .ZN(
        n23641) );
  OAI22_X2 U7877 ( .A1(n26371), .A2(n26797), .B1(n25814), .B2(n15628), .ZN(
        n23642) );
  OAI22_X2 U7879 ( .A1(n26371), .A2(n26798), .B1(n25811), .B2(n15628), .ZN(
        n23643) );
  OAI22_X2 U7881 ( .A1(n26371), .A2(n26799), .B1(n25808), .B2(n15628), .ZN(
        n23644) );
  OAI22_X2 U7883 ( .A1(n26371), .A2(n26800), .B1(n25805), .B2(n15628), .ZN(
        n23645) );
  OAI22_X2 U7885 ( .A1(n26371), .A2(n26801), .B1(n25802), .B2(n15628), .ZN(
        n23646) );
  OAI22_X2 U7887 ( .A1(n26371), .A2(n26802), .B1(n25797), .B2(n15628), .ZN(
        n23647) );
  OAI22_X2 U7889 ( .A1(n26371), .A2(n26803), .B1(n25792), .B2(n15628), .ZN(
        n23648) );
  OAI22_X2 U7891 ( .A1(n26371), .A2(n26804), .B1(n25790), .B2(n15628), .ZN(
        n23649) );
  OAI22_X2 U7893 ( .A1(n26371), .A2(n26805), .B1(n25787), .B2(n15628), .ZN(
        n23650) );
  OAI22_X2 U7895 ( .A1(n26371), .A2(n26806), .B1(n25784), .B2(n15628), .ZN(
        n23651) );
  OAI22_X2 U7899 ( .A1(n26370), .A2(n27047), .B1(n25834), .B2(n15631), .ZN(
        n23652) );
  OAI22_X2 U7901 ( .A1(n26370), .A2(n27048), .B1(n25828), .B2(n15631), .ZN(
        n23653) );
  OAI22_X2 U7903 ( .A1(n26370), .A2(n27049), .B1(n25826), .B2(n15631), .ZN(
        n23654) );
  OAI22_X2 U7905 ( .A1(n26370), .A2(n27050), .B1(n25823), .B2(n15631), .ZN(
        n23655) );
  OAI22_X2 U7907 ( .A1(n26370), .A2(n27051), .B1(n25820), .B2(n15631), .ZN(
        n23656) );
  OAI22_X2 U7909 ( .A1(n26370), .A2(n27052), .B1(n25817), .B2(n15631), .ZN(
        n23657) );
  OAI22_X2 U7911 ( .A1(n26370), .A2(n27053), .B1(n25814), .B2(n15631), .ZN(
        n23658) );
  OAI22_X2 U7913 ( .A1(n26370), .A2(n27054), .B1(n25811), .B2(n15631), .ZN(
        n23659) );
  OAI22_X2 U7915 ( .A1(n26370), .A2(n27055), .B1(n25808), .B2(n15631), .ZN(
        n23660) );
  OAI22_X2 U7917 ( .A1(n26370), .A2(n27056), .B1(n25805), .B2(n15631), .ZN(
        n23661) );
  OAI22_X2 U7919 ( .A1(n26370), .A2(n27057), .B1(n25802), .B2(n15631), .ZN(
        n23662) );
  OAI22_X2 U7921 ( .A1(n26370), .A2(n27058), .B1(n25797), .B2(n15631), .ZN(
        n23663) );
  OAI22_X2 U7923 ( .A1(n26370), .A2(n27059), .B1(n25792), .B2(n15631), .ZN(
        n23664) );
  OAI22_X2 U7925 ( .A1(n26370), .A2(n27060), .B1(n25790), .B2(n15631), .ZN(
        n23665) );
  OAI22_X2 U7927 ( .A1(n26370), .A2(n27061), .B1(n25787), .B2(n15631), .ZN(
        n23666) );
  OAI22_X2 U7929 ( .A1(n26370), .A2(n27062), .B1(n25784), .B2(n15631), .ZN(
        n23667) );
  OAI22_X2 U7933 ( .A1(n26369), .A2(n27303), .B1(n25832), .B2(n15649), .ZN(
        n23668) );
  OAI22_X2 U7935 ( .A1(n26369), .A2(n27304), .B1(n25828), .B2(n15649), .ZN(
        n23669) );
  OAI22_X2 U7937 ( .A1(n26369), .A2(n27305), .B1(n25824), .B2(n15649), .ZN(
        n23670) );
  OAI22_X2 U7939 ( .A1(n26369), .A2(n27306), .B1(n25821), .B2(n15649), .ZN(
        n23671) );
  OAI22_X2 U7941 ( .A1(n26369), .A2(n27307), .B1(n25818), .B2(n15649), .ZN(
        n23672) );
  OAI22_X2 U7943 ( .A1(n26369), .A2(n27308), .B1(n25815), .B2(n15649), .ZN(
        n23673) );
  OAI22_X2 U7945 ( .A1(n26369), .A2(n27309), .B1(n25812), .B2(n15649), .ZN(
        n23674) );
  OAI22_X2 U7947 ( .A1(n26369), .A2(n27310), .B1(n25809), .B2(n15649), .ZN(
        n23675) );
  OAI22_X2 U7949 ( .A1(n26369), .A2(n27311), .B1(n25806), .B2(n15649), .ZN(
        n23676) );
  OAI22_X2 U7951 ( .A1(n26369), .A2(n27312), .B1(n25803), .B2(n15649), .ZN(
        n23677) );
  OAI22_X2 U7953 ( .A1(n26369), .A2(n27313), .B1(n25800), .B2(n15649), .ZN(
        n23678) );
  OAI22_X2 U7955 ( .A1(n26369), .A2(n27314), .B1(n25797), .B2(n15649), .ZN(
        n23679) );
  OAI22_X2 U7957 ( .A1(n26369), .A2(n27315), .B1(n25792), .B2(n15649), .ZN(
        n23680) );
  OAI22_X2 U7959 ( .A1(n26369), .A2(n27316), .B1(n25788), .B2(n15649), .ZN(
        n23681) );
  OAI22_X2 U7961 ( .A1(n26369), .A2(n27317), .B1(n25785), .B2(n15649), .ZN(
        n23682) );
  OAI22_X2 U7963 ( .A1(n26369), .A2(n27318), .B1(n25782), .B2(n15649), .ZN(
        n23683) );
  OAI22_X2 U7968 ( .A1(n26364), .A2(n26647), .B1(n25833), .B2(n15667), .ZN(
        n23684) );
  OAI22_X2 U7970 ( .A1(n26364), .A2(n26648), .B1(n25828), .B2(n15667), .ZN(
        n23685) );
  OAI22_X2 U7972 ( .A1(n26364), .A2(n26649), .B1(n25825), .B2(n15667), .ZN(
        n23686) );
  OAI22_X2 U7974 ( .A1(n26364), .A2(n26650), .B1(n25822), .B2(n15667), .ZN(
        n23687) );
  OAI22_X2 U7976 ( .A1(n26364), .A2(n26651), .B1(n25819), .B2(n15667), .ZN(
        n23688) );
  OAI22_X2 U7978 ( .A1(n26364), .A2(n26652), .B1(n25816), .B2(n15667), .ZN(
        n23689) );
  OAI22_X2 U7980 ( .A1(n26364), .A2(n26653), .B1(n25813), .B2(n15667), .ZN(
        n23690) );
  OAI22_X2 U7982 ( .A1(n26364), .A2(n26654), .B1(n25810), .B2(n15667), .ZN(
        n23691) );
  OAI22_X2 U7984 ( .A1(n26364), .A2(n26655), .B1(n25807), .B2(n15667), .ZN(
        n23692) );
  OAI22_X2 U7986 ( .A1(n26364), .A2(n26656), .B1(n25804), .B2(n15667), .ZN(
        n23693) );
  OAI22_X2 U7988 ( .A1(n26364), .A2(n26657), .B1(n25801), .B2(n15667), .ZN(
        n23694) );
  OAI22_X2 U7990 ( .A1(n26364), .A2(n26658), .B1(n25797), .B2(n15667), .ZN(
        n23695) );
  OAI22_X2 U7992 ( .A1(n26364), .A2(n26659), .B1(n25792), .B2(n15667), .ZN(
        n23696) );
  OAI22_X2 U7994 ( .A1(n26364), .A2(n26660), .B1(n25789), .B2(n15667), .ZN(
        n23697) );
  OAI22_X2 U7996 ( .A1(n26364), .A2(n26661), .B1(n25786), .B2(n15667), .ZN(
        n23698) );
  OAI22_X2 U7998 ( .A1(n26364), .A2(n26662), .B1(n25783), .B2(n15667), .ZN(
        n23699) );
  OAI22_X2 U8002 ( .A1(n26363), .A2(n27575), .B1(n25832), .B2(n15684), .ZN(
        n23700) );
  OAI22_X2 U8004 ( .A1(n26363), .A2(n27576), .B1(n25828), .B2(n15684), .ZN(
        n23701) );
  OAI22_X2 U8006 ( .A1(n26363), .A2(n27577), .B1(n25824), .B2(n15684), .ZN(
        n23702) );
  OAI22_X2 U8008 ( .A1(n26363), .A2(n27578), .B1(n25821), .B2(n15684), .ZN(
        n23703) );
  OAI22_X2 U8010 ( .A1(n26363), .A2(n27579), .B1(n25818), .B2(n15684), .ZN(
        n23704) );
  OAI22_X2 U8012 ( .A1(n26363), .A2(n27580), .B1(n25815), .B2(n15684), .ZN(
        n23705) );
  OAI22_X2 U8014 ( .A1(n26363), .A2(n27581), .B1(n25812), .B2(n15684), .ZN(
        n23706) );
  OAI22_X2 U8016 ( .A1(n26363), .A2(n27582), .B1(n25809), .B2(n15684), .ZN(
        n23707) );
  OAI22_X2 U8018 ( .A1(n26363), .A2(n27583), .B1(n25806), .B2(n15684), .ZN(
        n23708) );
  OAI22_X2 U8020 ( .A1(n26363), .A2(n27584), .B1(n25803), .B2(n15684), .ZN(
        n23709) );
  OAI22_X2 U8022 ( .A1(n26363), .A2(n27585), .B1(n25800), .B2(n15684), .ZN(
        n23710) );
  OAI22_X2 U8024 ( .A1(n26363), .A2(n27586), .B1(n25797), .B2(n15684), .ZN(
        n23711) );
  OAI22_X2 U8026 ( .A1(n26363), .A2(n27587), .B1(n25792), .B2(n15684), .ZN(
        n23712) );
  OAI22_X2 U8028 ( .A1(n26363), .A2(n27588), .B1(n25788), .B2(n15684), .ZN(
        n23713) );
  OAI22_X2 U8030 ( .A1(n26363), .A2(n27589), .B1(n25785), .B2(n15684), .ZN(
        n23714) );
  OAI22_X2 U8032 ( .A1(n26363), .A2(n27590), .B1(n25782), .B2(n15684), .ZN(
        n23715) );
  OAI22_X2 U8036 ( .A1(n26362), .A2(n26807), .B1(n25833), .B2(n15686), .ZN(
        n23716) );
  OAI22_X2 U8038 ( .A1(n26362), .A2(n26808), .B1(n25828), .B2(n15686), .ZN(
        n23717) );
  OAI22_X2 U8040 ( .A1(n26362), .A2(n26809), .B1(n25825), .B2(n15686), .ZN(
        n23718) );
  OAI22_X2 U8042 ( .A1(n26362), .A2(n26810), .B1(n25822), .B2(n15686), .ZN(
        n23719) );
  OAI22_X2 U8044 ( .A1(n26362), .A2(n26811), .B1(n25819), .B2(n15686), .ZN(
        n23720) );
  OAI22_X2 U8046 ( .A1(n26362), .A2(n26812), .B1(n25816), .B2(n15686), .ZN(
        n23721) );
  OAI22_X2 U8048 ( .A1(n26362), .A2(n26813), .B1(n25813), .B2(n15686), .ZN(
        n23722) );
  OAI22_X2 U8050 ( .A1(n26362), .A2(n26814), .B1(n25810), .B2(n15686), .ZN(
        n23723) );
  OAI22_X2 U8052 ( .A1(n26362), .A2(n26815), .B1(n25807), .B2(n15686), .ZN(
        n23724) );
  OAI22_X2 U8054 ( .A1(n26362), .A2(n26816), .B1(n25804), .B2(n15686), .ZN(
        n23725) );
  OAI22_X2 U8056 ( .A1(n26362), .A2(n26817), .B1(n25801), .B2(n15686), .ZN(
        n23726) );
  OAI22_X2 U8058 ( .A1(n26362), .A2(n26818), .B1(n25797), .B2(n15686), .ZN(
        n23727) );
  OAI22_X2 U8060 ( .A1(n26362), .A2(n26819), .B1(n25792), .B2(n15686), .ZN(
        n23728) );
  OAI22_X2 U8062 ( .A1(n26362), .A2(n26820), .B1(n25789), .B2(n15686), .ZN(
        n23729) );
  OAI22_X2 U8064 ( .A1(n26362), .A2(n26821), .B1(n25786), .B2(n15686), .ZN(
        n23730) );
  OAI22_X2 U8066 ( .A1(n26362), .A2(n26822), .B1(n25783), .B2(n15686), .ZN(
        n23731) );
  OAI22_X2 U8070 ( .A1(n26361), .A2(n27063), .B1(n25834), .B2(n15689), .ZN(
        n23732) );
  OAI22_X2 U8072 ( .A1(n26361), .A2(n27064), .B1(n25828), .B2(n15689), .ZN(
        n23733) );
  OAI22_X2 U8074 ( .A1(n26361), .A2(n27065), .B1(n25826), .B2(n15689), .ZN(
        n23734) );
  OAI22_X2 U8076 ( .A1(n26361), .A2(n27066), .B1(n25823), .B2(n15689), .ZN(
        n23735) );
  OAI22_X2 U8078 ( .A1(n26361), .A2(n27067), .B1(n25820), .B2(n15689), .ZN(
        n23736) );
  OAI22_X2 U8080 ( .A1(n26361), .A2(n27068), .B1(n25817), .B2(n15689), .ZN(
        n23737) );
  OAI22_X2 U8082 ( .A1(n26361), .A2(n27069), .B1(n25814), .B2(n15689), .ZN(
        n23738) );
  OAI22_X2 U8084 ( .A1(n26361), .A2(n27070), .B1(n25811), .B2(n15689), .ZN(
        n23739) );
  OAI22_X2 U8086 ( .A1(n26361), .A2(n27071), .B1(n25808), .B2(n15689), .ZN(
        n23740) );
  OAI22_X2 U8088 ( .A1(n26361), .A2(n27072), .B1(n25805), .B2(n15689), .ZN(
        n23741) );
  OAI22_X2 U8090 ( .A1(n26361), .A2(n27073), .B1(n25802), .B2(n15689), .ZN(
        n23742) );
  OAI22_X2 U8092 ( .A1(n26361), .A2(n27074), .B1(n25797), .B2(n15689), .ZN(
        n23743) );
  OAI22_X2 U8094 ( .A1(n26361), .A2(n27075), .B1(n25792), .B2(n15689), .ZN(
        n23744) );
  OAI22_X2 U8096 ( .A1(n26361), .A2(n27076), .B1(n25790), .B2(n15689), .ZN(
        n23745) );
  OAI22_X2 U8098 ( .A1(n26361), .A2(n27077), .B1(n25787), .B2(n15689), .ZN(
        n23746) );
  OAI22_X2 U8100 ( .A1(n26361), .A2(n27078), .B1(n25784), .B2(n15689), .ZN(
        n23747) );
  OAI22_X2 U8104 ( .A1(n26360), .A2(n27319), .B1(n25833), .B2(n15707), .ZN(
        n23748) );
  OAI22_X2 U8106 ( .A1(n26360), .A2(n27320), .B1(n25829), .B2(n15707), .ZN(
        n23749) );
  OAI22_X2 U8108 ( .A1(n26360), .A2(n27321), .B1(n25825), .B2(n15707), .ZN(
        n23750) );
  OAI22_X2 U8110 ( .A1(n26360), .A2(n27322), .B1(n25822), .B2(n15707), .ZN(
        n23751) );
  OAI22_X2 U8112 ( .A1(n26360), .A2(n27323), .B1(n25819), .B2(n15707), .ZN(
        n23752) );
  OAI22_X2 U8114 ( .A1(n26360), .A2(n27324), .B1(n25816), .B2(n15707), .ZN(
        n23753) );
  OAI22_X2 U8116 ( .A1(n26360), .A2(n27325), .B1(n25813), .B2(n15707), .ZN(
        n23754) );
  OAI22_X2 U8118 ( .A1(n26360), .A2(n27326), .B1(n25810), .B2(n15707), .ZN(
        n23755) );
  OAI22_X2 U8120 ( .A1(n26360), .A2(n27327), .B1(n25807), .B2(n15707), .ZN(
        n23756) );
  OAI22_X2 U8122 ( .A1(n26360), .A2(n27328), .B1(n25804), .B2(n15707), .ZN(
        n23757) );
  OAI22_X2 U8124 ( .A1(n26360), .A2(n27329), .B1(n25801), .B2(n15707), .ZN(
        n23758) );
  OAI22_X2 U8126 ( .A1(n26360), .A2(n27330), .B1(n25798), .B2(n15707), .ZN(
        n23759) );
  OAI22_X2 U8128 ( .A1(n26360), .A2(n27331), .B1(n25793), .B2(n15707), .ZN(
        n23760) );
  OAI22_X2 U8130 ( .A1(n26360), .A2(n27332), .B1(n25789), .B2(n15707), .ZN(
        n23761) );
  OAI22_X2 U8132 ( .A1(n26360), .A2(n27333), .B1(n25786), .B2(n15707), .ZN(
        n23762) );
  OAI22_X2 U8134 ( .A1(n26360), .A2(n27334), .B1(n25783), .B2(n15707), .ZN(
        n23763) );
  OAI22_X2 U8139 ( .A1(n26355), .A2(n26567), .B1(n25833), .B2(n11430), .ZN(
        n23764) );
  OAI22_X2 U8141 ( .A1(n26355), .A2(n26568), .B1(n25831), .B2(n11430), .ZN(
        n23765) );
  OAI22_X2 U8143 ( .A1(n26355), .A2(n26569), .B1(n25825), .B2(n11430), .ZN(
        n23766) );
  OAI22_X2 U8145 ( .A1(n26355), .A2(n26570), .B1(n25822), .B2(n11430), .ZN(
        n23767) );
  OAI22_X2 U8147 ( .A1(n26355), .A2(n26571), .B1(n25819), .B2(n11430), .ZN(
        n23768) );
  OAI22_X2 U8149 ( .A1(n26355), .A2(n26572), .B1(n25816), .B2(n11430), .ZN(
        n23769) );
  OAI22_X2 U8151 ( .A1(n26355), .A2(n26573), .B1(n25813), .B2(n11430), .ZN(
        n23770) );
  OAI22_X2 U8153 ( .A1(n26355), .A2(n26574), .B1(n25810), .B2(n11430), .ZN(
        n23771) );
  OAI22_X2 U8155 ( .A1(n26355), .A2(n26575), .B1(n25807), .B2(n11430), .ZN(
        n23772) );
  OAI22_X2 U8157 ( .A1(n26355), .A2(n26576), .B1(n25804), .B2(n11430), .ZN(
        n23773) );
  OAI22_X2 U8159 ( .A1(n26355), .A2(n26577), .B1(n25801), .B2(n11430), .ZN(
        n23774) );
  OAI22_X2 U8161 ( .A1(n26355), .A2(n26578), .B1(n25798), .B2(n11430), .ZN(
        n23775) );
  OAI22_X2 U8163 ( .A1(n26355), .A2(n26579), .B1(n25795), .B2(n11430), .ZN(
        n23776) );
  OAI22_X2 U8165 ( .A1(n26355), .A2(n26580), .B1(n25789), .B2(n11430), .ZN(
        n23777) );
  OAI22_X2 U8167 ( .A1(n26355), .A2(n26581), .B1(n25786), .B2(n11430), .ZN(
        n23778) );
  OAI22_X2 U8169 ( .A1(n26355), .A2(n26582), .B1(n25783), .B2(n11430), .ZN(
        n23779) );
  OAI22_X2 U8173 ( .A1(n26354), .A2(n27591), .B1(n25833), .B2(n15741), .ZN(
        n23780) );
  OAI22_X2 U8175 ( .A1(n26354), .A2(n27592), .B1(n25829), .B2(n15741), .ZN(
        n23781) );
  OAI22_X2 U8177 ( .A1(n26354), .A2(n27593), .B1(n25825), .B2(n15741), .ZN(
        n23782) );
  OAI22_X2 U8179 ( .A1(n26354), .A2(n27594), .B1(n25822), .B2(n15741), .ZN(
        n23783) );
  OAI22_X2 U8181 ( .A1(n26354), .A2(n27595), .B1(n25819), .B2(n15741), .ZN(
        n23784) );
  OAI22_X2 U8183 ( .A1(n26354), .A2(n27596), .B1(n25816), .B2(n15741), .ZN(
        n23785) );
  OAI22_X2 U8185 ( .A1(n26354), .A2(n27597), .B1(n25813), .B2(n15741), .ZN(
        n23786) );
  OAI22_X2 U8187 ( .A1(n26354), .A2(n27598), .B1(n25810), .B2(n15741), .ZN(
        n23787) );
  OAI22_X2 U8189 ( .A1(n26354), .A2(n27599), .B1(n25807), .B2(n15741), .ZN(
        n23788) );
  OAI22_X2 U8191 ( .A1(n26354), .A2(n27600), .B1(n25804), .B2(n15741), .ZN(
        n23789) );
  OAI22_X2 U8193 ( .A1(n26354), .A2(n27601), .B1(n25801), .B2(n15741), .ZN(
        n23790) );
  OAI22_X2 U8195 ( .A1(n26354), .A2(n27602), .B1(n25798), .B2(n15741), .ZN(
        n23791) );
  OAI22_X2 U8197 ( .A1(n26354), .A2(n27603), .B1(n25793), .B2(n15741), .ZN(
        n23792) );
  OAI22_X2 U8199 ( .A1(n26354), .A2(n27604), .B1(n25789), .B2(n15741), .ZN(
        n23793) );
  OAI22_X2 U8201 ( .A1(n26354), .A2(n27605), .B1(n25786), .B2(n15741), .ZN(
        n23794) );
  OAI22_X2 U8203 ( .A1(n26354), .A2(n27606), .B1(n25783), .B2(n15741), .ZN(
        n23795) );
  OAI22_X2 U8207 ( .A1(n26353), .A2(n26823), .B1(n25832), .B2(n15743), .ZN(
        n23796) );
  OAI22_X2 U8209 ( .A1(n26353), .A2(n26824), .B1(n25829), .B2(n15743), .ZN(
        n23797) );
  OAI22_X2 U8211 ( .A1(n26353), .A2(n26825), .B1(n25824), .B2(n15743), .ZN(
        n23798) );
  OAI22_X2 U8213 ( .A1(n26353), .A2(n26826), .B1(n25821), .B2(n15743), .ZN(
        n23799) );
  OAI22_X2 U8215 ( .A1(n26353), .A2(n26827), .B1(n25818), .B2(n15743), .ZN(
        n23800) );
  OAI22_X2 U8217 ( .A1(n26353), .A2(n26828), .B1(n25815), .B2(n15743), .ZN(
        n23801) );
  OAI22_X2 U8219 ( .A1(n26353), .A2(n26829), .B1(n25812), .B2(n15743), .ZN(
        n23802) );
  OAI22_X2 U8221 ( .A1(n26353), .A2(n26830), .B1(n25809), .B2(n15743), .ZN(
        n23803) );
  OAI22_X2 U8223 ( .A1(n26353), .A2(n26831), .B1(n25806), .B2(n15743), .ZN(
        n23804) );
  OAI22_X2 U8225 ( .A1(n26353), .A2(n26832), .B1(n25803), .B2(n15743), .ZN(
        n23805) );
  OAI22_X2 U8227 ( .A1(n26353), .A2(n26833), .B1(n25800), .B2(n15743), .ZN(
        n23806) );
  OAI22_X2 U8229 ( .A1(n26353), .A2(n26834), .B1(n25798), .B2(n15743), .ZN(
        n23807) );
  OAI22_X2 U8231 ( .A1(n26353), .A2(n26835), .B1(n25793), .B2(n15743), .ZN(
        n23808) );
  OAI22_X2 U8233 ( .A1(n26353), .A2(n26836), .B1(n25788), .B2(n15743), .ZN(
        n23809) );
  OAI22_X2 U8235 ( .A1(n26353), .A2(n26837), .B1(n25785), .B2(n15743), .ZN(
        n23810) );
  OAI22_X2 U8237 ( .A1(n26353), .A2(n26838), .B1(n25782), .B2(n15743), .ZN(
        n23811) );
  OAI22_X2 U8241 ( .A1(n26352), .A2(n27079), .B1(n25834), .B2(n15746), .ZN(
        n23812) );
  OAI22_X2 U8243 ( .A1(n26352), .A2(n27080), .B1(n25829), .B2(n15746), .ZN(
        n23813) );
  OAI22_X2 U8245 ( .A1(n26352), .A2(n27081), .B1(n25826), .B2(n15746), .ZN(
        n23814) );
  OAI22_X2 U8247 ( .A1(n26352), .A2(n27082), .B1(n25823), .B2(n15746), .ZN(
        n23815) );
  OAI22_X2 U8249 ( .A1(n26352), .A2(n27083), .B1(n25820), .B2(n15746), .ZN(
        n23816) );
  OAI22_X2 U8251 ( .A1(n26352), .A2(n27084), .B1(n25817), .B2(n15746), .ZN(
        n23817) );
  OAI22_X2 U8253 ( .A1(n26352), .A2(n27085), .B1(n25814), .B2(n15746), .ZN(
        n23818) );
  OAI22_X2 U8255 ( .A1(n26352), .A2(n27086), .B1(n25811), .B2(n15746), .ZN(
        n23819) );
  OAI22_X2 U8257 ( .A1(n26352), .A2(n27087), .B1(n25808), .B2(n15746), .ZN(
        n23820) );
  OAI22_X2 U8259 ( .A1(n26352), .A2(n27088), .B1(n25805), .B2(n15746), .ZN(
        n23821) );
  OAI22_X2 U8261 ( .A1(n26352), .A2(n27089), .B1(n25802), .B2(n15746), .ZN(
        n23822) );
  OAI22_X2 U8263 ( .A1(n26352), .A2(n27090), .B1(n25798), .B2(n15746), .ZN(
        n23823) );
  OAI22_X2 U8265 ( .A1(n26352), .A2(n27091), .B1(n25793), .B2(n15746), .ZN(
        n23824) );
  OAI22_X2 U8267 ( .A1(n26352), .A2(n27092), .B1(n25790), .B2(n15746), .ZN(
        n23825) );
  OAI22_X2 U8269 ( .A1(n26352), .A2(n27093), .B1(n25787), .B2(n15746), .ZN(
        n23826) );
  OAI22_X2 U8271 ( .A1(n26352), .A2(n27094), .B1(n25784), .B2(n15746), .ZN(
        n23827) );
  OAI22_X2 U8275 ( .A1(n26351), .A2(n27335), .B1(n25833), .B2(n15764), .ZN(
        n23828) );
  OAI22_X2 U8277 ( .A1(n26351), .A2(n27336), .B1(n25829), .B2(n15764), .ZN(
        n23829) );
  OAI22_X2 U8279 ( .A1(n26351), .A2(n27337), .B1(n25825), .B2(n15764), .ZN(
        n23830) );
  OAI22_X2 U8281 ( .A1(n26351), .A2(n27338), .B1(n25822), .B2(n15764), .ZN(
        n23831) );
  OAI22_X2 U8283 ( .A1(n26351), .A2(n27339), .B1(n25819), .B2(n15764), .ZN(
        n23832) );
  OAI22_X2 U8285 ( .A1(n26351), .A2(n27340), .B1(n25816), .B2(n15764), .ZN(
        n23833) );
  OAI22_X2 U8287 ( .A1(n26351), .A2(n27341), .B1(n25813), .B2(n15764), .ZN(
        n23834) );
  OAI22_X2 U8289 ( .A1(n26351), .A2(n27342), .B1(n25810), .B2(n15764), .ZN(
        n23835) );
  OAI22_X2 U8291 ( .A1(n26351), .A2(n27343), .B1(n25807), .B2(n15764), .ZN(
        n23836) );
  OAI22_X2 U8293 ( .A1(n26351), .A2(n27344), .B1(n25804), .B2(n15764), .ZN(
        n23837) );
  OAI22_X2 U8295 ( .A1(n26351), .A2(n27345), .B1(n25801), .B2(n15764), .ZN(
        n23838) );
  OAI22_X2 U8297 ( .A1(n26351), .A2(n27346), .B1(n25798), .B2(n15764), .ZN(
        n23839) );
  OAI22_X2 U8299 ( .A1(n26351), .A2(n27347), .B1(n25793), .B2(n15764), .ZN(
        n23840) );
  OAI22_X2 U8301 ( .A1(n26351), .A2(n27348), .B1(n25789), .B2(n15764), .ZN(
        n23841) );
  OAI22_X2 U8303 ( .A1(n26351), .A2(n27349), .B1(n25786), .B2(n15764), .ZN(
        n23842) );
  OAI22_X2 U8305 ( .A1(n26351), .A2(n27350), .B1(n25783), .B2(n15764), .ZN(
        n23843) );
  NOR2_X2 U8310 ( .A1(n15780), .A2(n22381), .ZN(n15606) );
  OAI22_X2 U8311 ( .A1(n26418), .A2(n26519), .B1(n25832), .B2(n15782), .ZN(
        n23844) );
  OAI22_X2 U8313 ( .A1(n26418), .A2(n26520), .B1(n25829), .B2(n15782), .ZN(
        n23845) );
  OAI22_X2 U8315 ( .A1(n26418), .A2(n26521), .B1(n25824), .B2(n15782), .ZN(
        n23846) );
  OAI22_X2 U8317 ( .A1(n26418), .A2(n26522), .B1(n25821), .B2(n15782), .ZN(
        n23847) );
  OAI22_X2 U8319 ( .A1(n26418), .A2(n26523), .B1(n25818), .B2(n15782), .ZN(
        n23848) );
  OAI22_X2 U8321 ( .A1(n26418), .A2(n26524), .B1(n25815), .B2(n15782), .ZN(
        n23849) );
  OAI22_X2 U8323 ( .A1(n26418), .A2(n26525), .B1(n25812), .B2(n15782), .ZN(
        n23850) );
  OAI22_X2 U8325 ( .A1(n26418), .A2(n26526), .B1(n25809), .B2(n15782), .ZN(
        n23851) );
  OAI22_X2 U8327 ( .A1(n26418), .A2(n26527), .B1(n25806), .B2(n15782), .ZN(
        n23852) );
  OAI22_X2 U8329 ( .A1(n26418), .A2(n26528), .B1(n25803), .B2(n15782), .ZN(
        n23853) );
  OAI22_X2 U8331 ( .A1(n26418), .A2(n26529), .B1(n25800), .B2(n15782), .ZN(
        n23854) );
  OAI22_X2 U8333 ( .A1(n26418), .A2(n26530), .B1(n25798), .B2(n15782), .ZN(
        n23855) );
  OAI22_X2 U8335 ( .A1(n26418), .A2(n26531), .B1(n25793), .B2(n15782), .ZN(
        n23856) );
  OAI22_X2 U8337 ( .A1(n26418), .A2(n26532), .B1(n25788), .B2(n15782), .ZN(
        n23857) );
  OAI22_X2 U8339 ( .A1(n26418), .A2(n26533), .B1(n25785), .B2(n15782), .ZN(
        n23858) );
  OAI22_X2 U8341 ( .A1(n26418), .A2(n26534), .B1(n25782), .B2(n15782), .ZN(
        n23859) );
  OAI22_X2 U8345 ( .A1(n26417), .A2(n27607), .B1(n25832), .B2(n15785), .ZN(
        n23860) );
  OAI22_X2 U8347 ( .A1(n26417), .A2(n27608), .B1(n25829), .B2(n15785), .ZN(
        n23861) );
  OAI22_X2 U8349 ( .A1(n26417), .A2(n27609), .B1(n25824), .B2(n15785), .ZN(
        n23862) );
  OAI22_X2 U8351 ( .A1(n26417), .A2(n27610), .B1(n25821), .B2(n15785), .ZN(
        n23863) );
  OAI22_X2 U8353 ( .A1(n26417), .A2(n27611), .B1(n25818), .B2(n15785), .ZN(
        n23864) );
  OAI22_X2 U8355 ( .A1(n26417), .A2(n27612), .B1(n25815), .B2(n15785), .ZN(
        n23865) );
  OAI22_X2 U8357 ( .A1(n26417), .A2(n27613), .B1(n25812), .B2(n15785), .ZN(
        n23866) );
  OAI22_X2 U8359 ( .A1(n26417), .A2(n27614), .B1(n25809), .B2(n15785), .ZN(
        n23867) );
  OAI22_X2 U8361 ( .A1(n26417), .A2(n27615), .B1(n25806), .B2(n15785), .ZN(
        n23868) );
  OAI22_X2 U8363 ( .A1(n26417), .A2(n27616), .B1(n25803), .B2(n15785), .ZN(
        n23869) );
  OAI22_X2 U8365 ( .A1(n26417), .A2(n27617), .B1(n25800), .B2(n15785), .ZN(
        n23870) );
  OAI22_X2 U8367 ( .A1(n26417), .A2(n27618), .B1(n25798), .B2(n15785), .ZN(
        n23871) );
  OAI22_X2 U8369 ( .A1(n26417), .A2(n27619), .B1(n25793), .B2(n15785), .ZN(
        n23872) );
  OAI22_X2 U8371 ( .A1(n26417), .A2(n27620), .B1(n25788), .B2(n15785), .ZN(
        n23873) );
  OAI22_X2 U8373 ( .A1(n26417), .A2(n27621), .B1(n25785), .B2(n15785), .ZN(
        n23874) );
  OAI22_X2 U8375 ( .A1(n26417), .A2(n27622), .B1(n25782), .B2(n15785), .ZN(
        n23875) );
  OAI22_X2 U8379 ( .A1(n26416), .A2(n26839), .B1(n25834), .B2(n15803), .ZN(
        n23876) );
  OAI22_X2 U8381 ( .A1(n26416), .A2(n26840), .B1(n25829), .B2(n15803), .ZN(
        n23877) );
  OAI22_X2 U8383 ( .A1(n26416), .A2(n26841), .B1(n25826), .B2(n15803), .ZN(
        n23878) );
  OAI22_X2 U8385 ( .A1(n26416), .A2(n26842), .B1(n25823), .B2(n15803), .ZN(
        n23879) );
  OAI22_X2 U8387 ( .A1(n26416), .A2(n26843), .B1(n25820), .B2(n15803), .ZN(
        n23880) );
  OAI22_X2 U8389 ( .A1(n26416), .A2(n26844), .B1(n25817), .B2(n15803), .ZN(
        n23881) );
  OAI22_X2 U8391 ( .A1(n26416), .A2(n26845), .B1(n25814), .B2(n15803), .ZN(
        n23882) );
  OAI22_X2 U8393 ( .A1(n26416), .A2(n26846), .B1(n25811), .B2(n15803), .ZN(
        n23883) );
  OAI22_X2 U8395 ( .A1(n26416), .A2(n26847), .B1(n25808), .B2(n15803), .ZN(
        n23884) );
  OAI22_X2 U8397 ( .A1(n26416), .A2(n26848), .B1(n25805), .B2(n15803), .ZN(
        n23885) );
  OAI22_X2 U8399 ( .A1(n26416), .A2(n26849), .B1(n25802), .B2(n15803), .ZN(
        n23886) );
  OAI22_X2 U8401 ( .A1(n26416), .A2(n26850), .B1(n25798), .B2(n15803), .ZN(
        n23887) );
  OAI22_X2 U8403 ( .A1(n26416), .A2(n26851), .B1(n25793), .B2(n15803), .ZN(
        n23888) );
  OAI22_X2 U8405 ( .A1(n26416), .A2(n26852), .B1(n25790), .B2(n15803), .ZN(
        n23889) );
  OAI22_X2 U8407 ( .A1(n26416), .A2(n26853), .B1(n25787), .B2(n15803), .ZN(
        n23890) );
  OAI22_X2 U8409 ( .A1(n26416), .A2(n26854), .B1(n25784), .B2(n15803), .ZN(
        n23891) );
  OAI22_X2 U8413 ( .A1(n26415), .A2(n27095), .B1(n25833), .B2(n15820), .ZN(
        n23892) );
  OAI22_X2 U8415 ( .A1(n26415), .A2(n27096), .B1(n25829), .B2(n15820), .ZN(
        n23893) );
  OAI22_X2 U8417 ( .A1(n26415), .A2(n27097), .B1(n25825), .B2(n15820), .ZN(
        n23894) );
  OAI22_X2 U8419 ( .A1(n26415), .A2(n27098), .B1(n25822), .B2(n15820), .ZN(
        n23895) );
  OAI22_X2 U8421 ( .A1(n26415), .A2(n27099), .B1(n25819), .B2(n15820), .ZN(
        n23896) );
  OAI22_X2 U8423 ( .A1(n26415), .A2(n27100), .B1(n25816), .B2(n15820), .ZN(
        n23897) );
  OAI22_X2 U8425 ( .A1(n26415), .A2(n27101), .B1(n25813), .B2(n15820), .ZN(
        n23898) );
  OAI22_X2 U8427 ( .A1(n26415), .A2(n27102), .B1(n25810), .B2(n15820), .ZN(
        n23899) );
  OAI22_X2 U8429 ( .A1(n26415), .A2(n27103), .B1(n25807), .B2(n15820), .ZN(
        n23900) );
  OAI22_X2 U8431 ( .A1(n26415), .A2(n27104), .B1(n25804), .B2(n15820), .ZN(
        n23901) );
  OAI22_X2 U8433 ( .A1(n26415), .A2(n27105), .B1(n25801), .B2(n15820), .ZN(
        n23902) );
  OAI22_X2 U8435 ( .A1(n26415), .A2(n27106), .B1(n25798), .B2(n15820), .ZN(
        n23903) );
  OAI22_X2 U8437 ( .A1(n26415), .A2(n27107), .B1(n25793), .B2(n15820), .ZN(
        n23904) );
  OAI22_X2 U8439 ( .A1(n26415), .A2(n27108), .B1(n25789), .B2(n15820), .ZN(
        n23905) );
  OAI22_X2 U8441 ( .A1(n26415), .A2(n27109), .B1(n25786), .B2(n15820), .ZN(
        n23906) );
  OAI22_X2 U8443 ( .A1(n26415), .A2(n27110), .B1(n25783), .B2(n15820), .ZN(
        n23907) );
  OAI22_X2 U8447 ( .A1(n26414), .A2(n27351), .B1(n25832), .B2(n15822), .ZN(
        n23908) );
  OAI22_X2 U8449 ( .A1(n26414), .A2(n27352), .B1(n25829), .B2(n15822), .ZN(
        n23909) );
  OAI22_X2 U8451 ( .A1(n26414), .A2(n27353), .B1(n25824), .B2(n15822), .ZN(
        n23910) );
  OAI22_X2 U8453 ( .A1(n26414), .A2(n27354), .B1(n25821), .B2(n15822), .ZN(
        n23911) );
  OAI22_X2 U8455 ( .A1(n26414), .A2(n27355), .B1(n25818), .B2(n15822), .ZN(
        n23912) );
  OAI22_X2 U8457 ( .A1(n26414), .A2(n27356), .B1(n25815), .B2(n15822), .ZN(
        n23913) );
  OAI22_X2 U8459 ( .A1(n26414), .A2(n27357), .B1(n25812), .B2(n15822), .ZN(
        n23914) );
  OAI22_X2 U8461 ( .A1(n26414), .A2(n27358), .B1(n25809), .B2(n15822), .ZN(
        n23915) );
  OAI22_X2 U8463 ( .A1(n26414), .A2(n27359), .B1(n25806), .B2(n15822), .ZN(
        n23916) );
  OAI22_X2 U8465 ( .A1(n26414), .A2(n27360), .B1(n25803), .B2(n15822), .ZN(
        n23917) );
  OAI22_X2 U8467 ( .A1(n26414), .A2(n27361), .B1(n25800), .B2(n15822), .ZN(
        n23918) );
  OAI22_X2 U8469 ( .A1(n26414), .A2(n27362), .B1(n25798), .B2(n15822), .ZN(
        n23919) );
  OAI22_X2 U8471 ( .A1(n26414), .A2(n27363), .B1(n25793), .B2(n15822), .ZN(
        n23920) );
  OAI22_X2 U8473 ( .A1(n26414), .A2(n27364), .B1(n25788), .B2(n15822), .ZN(
        n23921) );
  OAI22_X2 U8475 ( .A1(n26414), .A2(n27365), .B1(n25785), .B2(n15822), .ZN(
        n23922) );
  OAI22_X2 U8477 ( .A1(n26414), .A2(n27366), .B1(n25782), .B2(n15822), .ZN(
        n23923) );
  OAI22_X2 U8482 ( .A1(n26409), .A2(n26727), .B1(n25834), .B2(n15825), .ZN(
        n23924) );
  OAI22_X2 U8484 ( .A1(n26409), .A2(n26728), .B1(n25829), .B2(n15825), .ZN(
        n23925) );
  OAI22_X2 U8486 ( .A1(n26409), .A2(n26729), .B1(n25826), .B2(n15825), .ZN(
        n23926) );
  OAI22_X2 U8488 ( .A1(n26409), .A2(n26730), .B1(n25823), .B2(n15825), .ZN(
        n23927) );
  OAI22_X2 U8490 ( .A1(n26409), .A2(n26731), .B1(n25820), .B2(n15825), .ZN(
        n23928) );
  OAI22_X2 U8492 ( .A1(n26409), .A2(n26732), .B1(n25817), .B2(n15825), .ZN(
        n23929) );
  OAI22_X2 U8494 ( .A1(n26409), .A2(n26733), .B1(n25814), .B2(n15825), .ZN(
        n23930) );
  OAI22_X2 U8496 ( .A1(n26409), .A2(n26734), .B1(n25811), .B2(n15825), .ZN(
        n23931) );
  OAI22_X2 U8498 ( .A1(n26409), .A2(n26735), .B1(n25808), .B2(n15825), .ZN(
        n23932) );
  OAI22_X2 U8500 ( .A1(n26409), .A2(n26736), .B1(n25805), .B2(n15825), .ZN(
        n23933) );
  OAI22_X2 U8502 ( .A1(n26409), .A2(n26737), .B1(n25802), .B2(n15825), .ZN(
        n23934) );
  OAI22_X2 U8504 ( .A1(n26409), .A2(n26738), .B1(n25798), .B2(n15825), .ZN(
        n23935) );
  OAI22_X2 U8506 ( .A1(n26409), .A2(n26739), .B1(n25793), .B2(n15825), .ZN(
        n23936) );
  OAI22_X2 U8508 ( .A1(n26409), .A2(n26740), .B1(n25790), .B2(n15825), .ZN(
        n23937) );
  OAI22_X2 U8510 ( .A1(n26409), .A2(n26741), .B1(n25787), .B2(n15825), .ZN(
        n23938) );
  OAI22_X2 U8512 ( .A1(n26409), .A2(n26742), .B1(n25784), .B2(n15825), .ZN(
        n23939) );
  OAI22_X2 U8516 ( .A1(n26408), .A2(n27623), .B1(n25834), .B2(n15828), .ZN(
        n23940) );
  OAI22_X2 U8518 ( .A1(n26408), .A2(n27624), .B1(n25829), .B2(n15828), .ZN(
        n23941) );
  OAI22_X2 U8520 ( .A1(n26408), .A2(n27625), .B1(n25826), .B2(n15828), .ZN(
        n23942) );
  OAI22_X2 U8522 ( .A1(n26408), .A2(n27626), .B1(n25823), .B2(n15828), .ZN(
        n23943) );
  OAI22_X2 U8524 ( .A1(n26408), .A2(n27627), .B1(n25820), .B2(n15828), .ZN(
        n23944) );
  OAI22_X2 U8526 ( .A1(n26408), .A2(n27628), .B1(n25817), .B2(n15828), .ZN(
        n23945) );
  OAI22_X2 U8528 ( .A1(n26408), .A2(n27629), .B1(n25814), .B2(n15828), .ZN(
        n23946) );
  OAI22_X2 U8530 ( .A1(n26408), .A2(n27630), .B1(n25811), .B2(n15828), .ZN(
        n23947) );
  OAI22_X2 U8532 ( .A1(n26408), .A2(n27631), .B1(n25808), .B2(n15828), .ZN(
        n23948) );
  OAI22_X2 U8534 ( .A1(n26408), .A2(n27632), .B1(n25805), .B2(n15828), .ZN(
        n23949) );
  OAI22_X2 U8536 ( .A1(n26408), .A2(n27633), .B1(n25802), .B2(n15828), .ZN(
        n23950) );
  OAI22_X2 U8538 ( .A1(n26408), .A2(n27634), .B1(n25798), .B2(n15828), .ZN(
        n23951) );
  OAI22_X2 U8540 ( .A1(n26408), .A2(n27635), .B1(n25793), .B2(n15828), .ZN(
        n23952) );
  OAI22_X2 U8542 ( .A1(n26408), .A2(n27636), .B1(n25790), .B2(n15828), .ZN(
        n23953) );
  OAI22_X2 U8544 ( .A1(n26408), .A2(n27637), .B1(n25787), .B2(n15828), .ZN(
        n23954) );
  OAI22_X2 U8546 ( .A1(n26408), .A2(n27638), .B1(n25784), .B2(n15828), .ZN(
        n23955) );
  OAI22_X2 U8550 ( .A1(n26407), .A2(n26855), .B1(n25833), .B2(n15846), .ZN(
        n23956) );
  OAI22_X2 U8552 ( .A1(n26407), .A2(n26856), .B1(n25829), .B2(n15846), .ZN(
        n23957) );
  OAI22_X2 U8554 ( .A1(n26407), .A2(n26857), .B1(n25825), .B2(n15846), .ZN(
        n23958) );
  OAI22_X2 U8556 ( .A1(n26407), .A2(n26858), .B1(n25822), .B2(n15846), .ZN(
        n23959) );
  OAI22_X2 U8558 ( .A1(n26407), .A2(n26859), .B1(n25819), .B2(n15846), .ZN(
        n23960) );
  OAI22_X2 U8560 ( .A1(n26407), .A2(n26860), .B1(n25816), .B2(n15846), .ZN(
        n23961) );
  OAI22_X2 U8562 ( .A1(n26407), .A2(n26861), .B1(n25813), .B2(n15846), .ZN(
        n23962) );
  OAI22_X2 U8564 ( .A1(n26407), .A2(n26862), .B1(n25810), .B2(n15846), .ZN(
        n23963) );
  OAI22_X2 U8566 ( .A1(n26407), .A2(n26863), .B1(n25807), .B2(n15846), .ZN(
        n23964) );
  OAI22_X2 U8568 ( .A1(n26407), .A2(n26864), .B1(n25804), .B2(n15846), .ZN(
        n23965) );
  OAI22_X2 U8570 ( .A1(n26407), .A2(n26865), .B1(n25801), .B2(n15846), .ZN(
        n23966) );
  OAI22_X2 U8572 ( .A1(n26407), .A2(n26866), .B1(n25798), .B2(n15846), .ZN(
        n23967) );
  OAI22_X2 U8574 ( .A1(n26407), .A2(n26867), .B1(n25793), .B2(n15846), .ZN(
        n23968) );
  OAI22_X2 U8576 ( .A1(n26407), .A2(n26868), .B1(n25789), .B2(n15846), .ZN(
        n23969) );
  OAI22_X2 U8578 ( .A1(n26407), .A2(n26869), .B1(n25786), .B2(n15846), .ZN(
        n23970) );
  OAI22_X2 U8580 ( .A1(n26407), .A2(n26870), .B1(n25783), .B2(n15846), .ZN(
        n23971) );
  OAI22_X2 U8584 ( .A1(n26406), .A2(n27111), .B1(n25832), .B2(n15863), .ZN(
        n23972) );
  OAI22_X2 U8586 ( .A1(n26406), .A2(n27112), .B1(n25829), .B2(n15863), .ZN(
        n23973) );
  OAI22_X2 U8588 ( .A1(n26406), .A2(n27113), .B1(n25824), .B2(n15863), .ZN(
        n23974) );
  OAI22_X2 U8590 ( .A1(n26406), .A2(n27114), .B1(n25821), .B2(n15863), .ZN(
        n23975) );
  OAI22_X2 U8592 ( .A1(n26406), .A2(n27115), .B1(n25818), .B2(n15863), .ZN(
        n23976) );
  OAI22_X2 U8594 ( .A1(n26406), .A2(n27116), .B1(n25815), .B2(n15863), .ZN(
        n23977) );
  OAI22_X2 U8596 ( .A1(n26406), .A2(n27117), .B1(n25812), .B2(n15863), .ZN(
        n23978) );
  OAI22_X2 U8598 ( .A1(n26406), .A2(n27118), .B1(n25809), .B2(n15863), .ZN(
        n23979) );
  OAI22_X2 U8600 ( .A1(n26406), .A2(n27119), .B1(n25806), .B2(n15863), .ZN(
        n23980) );
  OAI22_X2 U8602 ( .A1(n26406), .A2(n27120), .B1(n25803), .B2(n15863), .ZN(
        n23981) );
  OAI22_X2 U8604 ( .A1(n26406), .A2(n27121), .B1(n25800), .B2(n15863), .ZN(
        n23982) );
  OAI22_X2 U8606 ( .A1(n26406), .A2(n27122), .B1(n25798), .B2(n15863), .ZN(
        n23983) );
  OAI22_X2 U8608 ( .A1(n26406), .A2(n27123), .B1(n25793), .B2(n15863), .ZN(
        n23984) );
  OAI22_X2 U8610 ( .A1(n26406), .A2(n27124), .B1(n25788), .B2(n15863), .ZN(
        n23985) );
  OAI22_X2 U8612 ( .A1(n26406), .A2(n27125), .B1(n25785), .B2(n15863), .ZN(
        n23986) );
  OAI22_X2 U8614 ( .A1(n26406), .A2(n27126), .B1(n25782), .B2(n15863), .ZN(
        n23987) );
  OAI22_X2 U8618 ( .A1(n26405), .A2(n27367), .B1(n25834), .B2(n15865), .ZN(
        n23988) );
  OAI22_X2 U8620 ( .A1(n26405), .A2(n27368), .B1(n25829), .B2(n15865), .ZN(
        n23989) );
  OAI22_X2 U8622 ( .A1(n26405), .A2(n27369), .B1(n25826), .B2(n15865), .ZN(
        n23990) );
  OAI22_X2 U8624 ( .A1(n26405), .A2(n27370), .B1(n25823), .B2(n15865), .ZN(
        n23991) );
  OAI22_X2 U8626 ( .A1(n26405), .A2(n27371), .B1(n25820), .B2(n15865), .ZN(
        n23992) );
  OAI22_X2 U8628 ( .A1(n26405), .A2(n27372), .B1(n25817), .B2(n15865), .ZN(
        n23993) );
  OAI22_X2 U8630 ( .A1(n26405), .A2(n27373), .B1(n25814), .B2(n15865), .ZN(
        n23994) );
  OAI22_X2 U8632 ( .A1(n26405), .A2(n27374), .B1(n25811), .B2(n15865), .ZN(
        n23995) );
  OAI22_X2 U8634 ( .A1(n26405), .A2(n27375), .B1(n25808), .B2(n15865), .ZN(
        n23996) );
  OAI22_X2 U8636 ( .A1(n26405), .A2(n27376), .B1(n25805), .B2(n15865), .ZN(
        n23997) );
  OAI22_X2 U8638 ( .A1(n26405), .A2(n27377), .B1(n25802), .B2(n15865), .ZN(
        n23998) );
  OAI22_X2 U8640 ( .A1(n26405), .A2(n27378), .B1(n25798), .B2(n15865), .ZN(
        n23999) );
  OAI22_X2 U8642 ( .A1(n26405), .A2(n27379), .B1(n25793), .B2(n15865), .ZN(
        n24000) );
  OAI22_X2 U8644 ( .A1(n26405), .A2(n27380), .B1(n25790), .B2(n15865), .ZN(
        n24001) );
  OAI22_X2 U8646 ( .A1(n26405), .A2(n27381), .B1(n25787), .B2(n15865), .ZN(
        n24002) );
  OAI22_X2 U8648 ( .A1(n26405), .A2(n27382), .B1(n25784), .B2(n15865), .ZN(
        n24003) );
  OAI22_X2 U8653 ( .A1(n26400), .A2(n26663), .B1(n25833), .B2(n15867), .ZN(
        n24004) );
  OAI22_X2 U8655 ( .A1(n26400), .A2(n26664), .B1(n25829), .B2(n15867), .ZN(
        n24005) );
  OAI22_X2 U8657 ( .A1(n26400), .A2(n26665), .B1(n25825), .B2(n15867), .ZN(
        n24006) );
  OAI22_X2 U8659 ( .A1(n26400), .A2(n26666), .B1(n25822), .B2(n15867), .ZN(
        n24007) );
  OAI22_X2 U8661 ( .A1(n26400), .A2(n26667), .B1(n25819), .B2(n15867), .ZN(
        n24008) );
  OAI22_X2 U8663 ( .A1(n26400), .A2(n26668), .B1(n25816), .B2(n15867), .ZN(
        n24009) );
  OAI22_X2 U8665 ( .A1(n26400), .A2(n26669), .B1(n25813), .B2(n15867), .ZN(
        n24010) );
  OAI22_X2 U8667 ( .A1(n26400), .A2(n26670), .B1(n25810), .B2(n15867), .ZN(
        n24011) );
  OAI22_X2 U8669 ( .A1(n26400), .A2(n26671), .B1(n25807), .B2(n15867), .ZN(
        n24012) );
  OAI22_X2 U8671 ( .A1(n26400), .A2(n26672), .B1(n25804), .B2(n15867), .ZN(
        n24013) );
  OAI22_X2 U8673 ( .A1(n26400), .A2(n26673), .B1(n25801), .B2(n15867), .ZN(
        n24014) );
  OAI22_X2 U8675 ( .A1(n26400), .A2(n26674), .B1(n25798), .B2(n15867), .ZN(
        n24015) );
  OAI22_X2 U8677 ( .A1(n26400), .A2(n26675), .B1(n25793), .B2(n15867), .ZN(
        n24016) );
  OAI22_X2 U8679 ( .A1(n26400), .A2(n26676), .B1(n25789), .B2(n15867), .ZN(
        n24017) );
  OAI22_X2 U8681 ( .A1(n26400), .A2(n26677), .B1(n25786), .B2(n15867), .ZN(
        n24018) );
  OAI22_X2 U8683 ( .A1(n26400), .A2(n26678), .B1(n25783), .B2(n15867), .ZN(
        n24019) );
  OAI22_X2 U8687 ( .A1(n26399), .A2(n27639), .B1(n25833), .B2(n15870), .ZN(
        n24020) );
  OAI22_X2 U8689 ( .A1(n26399), .A2(n27640), .B1(n25829), .B2(n15870), .ZN(
        n24021) );
  OAI22_X2 U8691 ( .A1(n26399), .A2(n27641), .B1(n25825), .B2(n15870), .ZN(
        n24022) );
  OAI22_X2 U8693 ( .A1(n26399), .A2(n27642), .B1(n25822), .B2(n15870), .ZN(
        n24023) );
  OAI22_X2 U8695 ( .A1(n26399), .A2(n27643), .B1(n25819), .B2(n15870), .ZN(
        n24024) );
  OAI22_X2 U8697 ( .A1(n26399), .A2(n27644), .B1(n25816), .B2(n15870), .ZN(
        n24025) );
  OAI22_X2 U8699 ( .A1(n26399), .A2(n27645), .B1(n25813), .B2(n15870), .ZN(
        n24026) );
  OAI22_X2 U8701 ( .A1(n26399), .A2(n27646), .B1(n25810), .B2(n15870), .ZN(
        n24027) );
  OAI22_X2 U8703 ( .A1(n26399), .A2(n27647), .B1(n25807), .B2(n15870), .ZN(
        n24028) );
  OAI22_X2 U8705 ( .A1(n26399), .A2(n27648), .B1(n25804), .B2(n15870), .ZN(
        n24029) );
  OAI22_X2 U8707 ( .A1(n26399), .A2(n27649), .B1(n25801), .B2(n15870), .ZN(
        n24030) );
  OAI22_X2 U8709 ( .A1(n26399), .A2(n27650), .B1(n25798), .B2(n15870), .ZN(
        n24031) );
  OAI22_X2 U8711 ( .A1(n26399), .A2(n27651), .B1(n25793), .B2(n15870), .ZN(
        n24032) );
  OAI22_X2 U8713 ( .A1(n26399), .A2(n27652), .B1(n25789), .B2(n15870), .ZN(
        n24033) );
  OAI22_X2 U8715 ( .A1(n26399), .A2(n27653), .B1(n25786), .B2(n15870), .ZN(
        n24034) );
  OAI22_X2 U8717 ( .A1(n26399), .A2(n27654), .B1(n25783), .B2(n15870), .ZN(
        n24035) );
  OAI22_X2 U8721 ( .A1(n26398), .A2(n26871), .B1(n25832), .B2(n15888), .ZN(
        n24036) );
  OAI22_X2 U8723 ( .A1(n26398), .A2(n26872), .B1(n25829), .B2(n15888), .ZN(
        n24037) );
  OAI22_X2 U8725 ( .A1(n26398), .A2(n26873), .B1(n25824), .B2(n15888), .ZN(
        n24038) );
  OAI22_X2 U8727 ( .A1(n26398), .A2(n26874), .B1(n25821), .B2(n15888), .ZN(
        n24039) );
  OAI22_X2 U8729 ( .A1(n26398), .A2(n26875), .B1(n25818), .B2(n15888), .ZN(
        n24040) );
  OAI22_X2 U8731 ( .A1(n26398), .A2(n26876), .B1(n25815), .B2(n15888), .ZN(
        n24041) );
  OAI22_X2 U8733 ( .A1(n26398), .A2(n26877), .B1(n25812), .B2(n15888), .ZN(
        n24042) );
  OAI22_X2 U8735 ( .A1(n26398), .A2(n26878), .B1(n25809), .B2(n15888), .ZN(
        n24043) );
  OAI22_X2 U8737 ( .A1(n26398), .A2(n26879), .B1(n25806), .B2(n15888), .ZN(
        n24044) );
  OAI22_X2 U8739 ( .A1(n26398), .A2(n26880), .B1(n25803), .B2(n15888), .ZN(
        n24045) );
  OAI22_X2 U8741 ( .A1(n26398), .A2(n26881), .B1(n25800), .B2(n15888), .ZN(
        n24046) );
  OAI22_X2 U8743 ( .A1(n26398), .A2(n26882), .B1(n25798), .B2(n15888), .ZN(
        n24047) );
  OAI22_X2 U8745 ( .A1(n26398), .A2(n26883), .B1(n25793), .B2(n15888), .ZN(
        n24048) );
  OAI22_X2 U8747 ( .A1(n26398), .A2(n26884), .B1(n25788), .B2(n15888), .ZN(
        n24049) );
  OAI22_X2 U8749 ( .A1(n26398), .A2(n26885), .B1(n25785), .B2(n15888), .ZN(
        n24050) );
  OAI22_X2 U8751 ( .A1(n26398), .A2(n26886), .B1(n25782), .B2(n15888), .ZN(
        n24051) );
  OAI22_X2 U8755 ( .A1(n26397), .A2(n27127), .B1(n25834), .B2(n15905), .ZN(
        n24052) );
  OAI22_X2 U8757 ( .A1(n26397), .A2(n27128), .B1(n25829), .B2(n15905), .ZN(
        n24053) );
  OAI22_X2 U8759 ( .A1(n26397), .A2(n27129), .B1(n25826), .B2(n15905), .ZN(
        n24054) );
  OAI22_X2 U8761 ( .A1(n26397), .A2(n27130), .B1(n25823), .B2(n15905), .ZN(
        n24055) );
  OAI22_X2 U8763 ( .A1(n26397), .A2(n27131), .B1(n25820), .B2(n15905), .ZN(
        n24056) );
  OAI22_X2 U8765 ( .A1(n26397), .A2(n27132), .B1(n25817), .B2(n15905), .ZN(
        n24057) );
  OAI22_X2 U8767 ( .A1(n26397), .A2(n27133), .B1(n25814), .B2(n15905), .ZN(
        n24058) );
  OAI22_X2 U8769 ( .A1(n26397), .A2(n27134), .B1(n25811), .B2(n15905), .ZN(
        n24059) );
  OAI22_X2 U8771 ( .A1(n26397), .A2(n27135), .B1(n25808), .B2(n15905), .ZN(
        n24060) );
  OAI22_X2 U8773 ( .A1(n26397), .A2(n27136), .B1(n25805), .B2(n15905), .ZN(
        n24061) );
  OAI22_X2 U8775 ( .A1(n26397), .A2(n27137), .B1(n25802), .B2(n15905), .ZN(
        n24062) );
  OAI22_X2 U8777 ( .A1(n26397), .A2(n27138), .B1(n25798), .B2(n15905), .ZN(
        n24063) );
  OAI22_X2 U8779 ( .A1(n26397), .A2(n27139), .B1(n25793), .B2(n15905), .ZN(
        n24064) );
  OAI22_X2 U8781 ( .A1(n26397), .A2(n27140), .B1(n25790), .B2(n15905), .ZN(
        n24065) );
  OAI22_X2 U8783 ( .A1(n26397), .A2(n27141), .B1(n25787), .B2(n15905), .ZN(
        n24066) );
  OAI22_X2 U8785 ( .A1(n26397), .A2(n27142), .B1(n25784), .B2(n15905), .ZN(
        n24067) );
  OAI22_X2 U8789 ( .A1(n26396), .A2(n27383), .B1(n25833), .B2(n15907), .ZN(
        n24068) );
  OAI22_X2 U8791 ( .A1(n26396), .A2(n27384), .B1(n25829), .B2(n15907), .ZN(
        n24069) );
  OAI22_X2 U8793 ( .A1(n26396), .A2(n27385), .B1(n25825), .B2(n15907), .ZN(
        n24070) );
  OAI22_X2 U8795 ( .A1(n26396), .A2(n27386), .B1(n25822), .B2(n15907), .ZN(
        n24071) );
  OAI22_X2 U8797 ( .A1(n26396), .A2(n27387), .B1(n25819), .B2(n15907), .ZN(
        n24072) );
  OAI22_X2 U8799 ( .A1(n26396), .A2(n27388), .B1(n25816), .B2(n15907), .ZN(
        n24073) );
  OAI22_X2 U8801 ( .A1(n26396), .A2(n27389), .B1(n25813), .B2(n15907), .ZN(
        n24074) );
  OAI22_X2 U8803 ( .A1(n26396), .A2(n27390), .B1(n25810), .B2(n15907), .ZN(
        n24075) );
  OAI22_X2 U8805 ( .A1(n26396), .A2(n27391), .B1(n25807), .B2(n15907), .ZN(
        n24076) );
  OAI22_X2 U8807 ( .A1(n26396), .A2(n27392), .B1(n25804), .B2(n15907), .ZN(
        n24077) );
  OAI22_X2 U8809 ( .A1(n26396), .A2(n27393), .B1(n25801), .B2(n15907), .ZN(
        n24078) );
  OAI22_X2 U8811 ( .A1(n26396), .A2(n27394), .B1(n25798), .B2(n15907), .ZN(
        n24079) );
  OAI22_X2 U8813 ( .A1(n26396), .A2(n27395), .B1(n25793), .B2(n15907), .ZN(
        n24080) );
  OAI22_X2 U8815 ( .A1(n26396), .A2(n27396), .B1(n25789), .B2(n15907), .ZN(
        n24081) );
  OAI22_X2 U8817 ( .A1(n26396), .A2(n27397), .B1(n25786), .B2(n15907), .ZN(
        n24082) );
  OAI22_X2 U8819 ( .A1(n26396), .A2(n27398), .B1(n25783), .B2(n15907), .ZN(
        n24083) );
  OAI22_X2 U8824 ( .A1(n26391), .A2(n26535), .B1(n25832), .B2(n15909), .ZN(
        n24084) );
  OAI22_X2 U8826 ( .A1(n26391), .A2(n26536), .B1(n25829), .B2(n15909), .ZN(
        n24085) );
  OAI22_X2 U8828 ( .A1(n26391), .A2(n26537), .B1(n25824), .B2(n15909), .ZN(
        n24086) );
  OAI22_X2 U8830 ( .A1(n26391), .A2(n26538), .B1(n25821), .B2(n15909), .ZN(
        n24087) );
  OAI22_X2 U8832 ( .A1(n26391), .A2(n26539), .B1(n25818), .B2(n15909), .ZN(
        n24088) );
  OAI22_X2 U8834 ( .A1(n26391), .A2(n26540), .B1(n25815), .B2(n15909), .ZN(
        n24089) );
  OAI22_X2 U8836 ( .A1(n26391), .A2(n26541), .B1(n25812), .B2(n15909), .ZN(
        n24090) );
  OAI22_X2 U8838 ( .A1(n26391), .A2(n26542), .B1(n25809), .B2(n15909), .ZN(
        n24091) );
  OAI22_X2 U8840 ( .A1(n26391), .A2(n26543), .B1(n25806), .B2(n15909), .ZN(
        n24092) );
  OAI22_X2 U8842 ( .A1(n26391), .A2(n26544), .B1(n25803), .B2(n15909), .ZN(
        n24093) );
  OAI22_X2 U8844 ( .A1(n26391), .A2(n26545), .B1(n25800), .B2(n15909), .ZN(
        n24094) );
  OAI22_X2 U8846 ( .A1(n26391), .A2(n26546), .B1(n25798), .B2(n15909), .ZN(
        n24095) );
  OAI22_X2 U8848 ( .A1(n26391), .A2(n26547), .B1(n25793), .B2(n15909), .ZN(
        n24096) );
  OAI22_X2 U8850 ( .A1(n26391), .A2(n26548), .B1(n25788), .B2(n15909), .ZN(
        n24097) );
  OAI22_X2 U8852 ( .A1(n26391), .A2(n26549), .B1(n25785), .B2(n15909), .ZN(
        n24098) );
  OAI22_X2 U8854 ( .A1(n26391), .A2(n26550), .B1(n25782), .B2(n15909), .ZN(
        n24099) );
  OAI22_X2 U8858 ( .A1(n26390), .A2(n27655), .B1(n25832), .B2(n15912), .ZN(
        n24100) );
  OAI22_X2 U8860 ( .A1(n26390), .A2(n27656), .B1(n25829), .B2(n15912), .ZN(
        n24101) );
  OAI22_X2 U8862 ( .A1(n26390), .A2(n27657), .B1(n25824), .B2(n15912), .ZN(
        n24102) );
  OAI22_X2 U8864 ( .A1(n26390), .A2(n27658), .B1(n25821), .B2(n15912), .ZN(
        n24103) );
  OAI22_X2 U8866 ( .A1(n26390), .A2(n27659), .B1(n25818), .B2(n15912), .ZN(
        n24104) );
  OAI22_X2 U8868 ( .A1(n26390), .A2(n27660), .B1(n25815), .B2(n15912), .ZN(
        n24105) );
  OAI22_X2 U8870 ( .A1(n26390), .A2(n27661), .B1(n25812), .B2(n15912), .ZN(
        n24106) );
  OAI22_X2 U8872 ( .A1(n26390), .A2(n27662), .B1(n25809), .B2(n15912), .ZN(
        n24107) );
  OAI22_X2 U8874 ( .A1(n26390), .A2(n27663), .B1(n25806), .B2(n15912), .ZN(
        n24108) );
  OAI22_X2 U8876 ( .A1(n26390), .A2(n27664), .B1(n25803), .B2(n15912), .ZN(
        n24109) );
  OAI22_X2 U8878 ( .A1(n26390), .A2(n27665), .B1(n25800), .B2(n15912), .ZN(
        n24110) );
  OAI22_X2 U8880 ( .A1(n26390), .A2(n27666), .B1(n25798), .B2(n15912), .ZN(
        n24111) );
  OAI22_X2 U8882 ( .A1(n26390), .A2(n27667), .B1(n25793), .B2(n15912), .ZN(
        n24112) );
  OAI22_X2 U8884 ( .A1(n26390), .A2(n27668), .B1(n25788), .B2(n15912), .ZN(
        n24113) );
  OAI22_X2 U8886 ( .A1(n26390), .A2(n27669), .B1(n25785), .B2(n15912), .ZN(
        n24114) );
  OAI22_X2 U8888 ( .A1(n26390), .A2(n27670), .B1(n25782), .B2(n15912), .ZN(
        n24115) );
  OAI22_X2 U8892 ( .A1(n26389), .A2(n26887), .B1(n25834), .B2(n15930), .ZN(
        n24116) );
  OAI22_X2 U8894 ( .A1(n26389), .A2(n26888), .B1(n25829), .B2(n15930), .ZN(
        n24117) );
  OAI22_X2 U8896 ( .A1(n26389), .A2(n26889), .B1(n25826), .B2(n15930), .ZN(
        n24118) );
  OAI22_X2 U8898 ( .A1(n26389), .A2(n26890), .B1(n25823), .B2(n15930), .ZN(
        n24119) );
  OAI22_X2 U8900 ( .A1(n26389), .A2(n26891), .B1(n25820), .B2(n15930), .ZN(
        n24120) );
  OAI22_X2 U8902 ( .A1(n26389), .A2(n26892), .B1(n25817), .B2(n15930), .ZN(
        n24121) );
  OAI22_X2 U8904 ( .A1(n26389), .A2(n26893), .B1(n25814), .B2(n15930), .ZN(
        n24122) );
  OAI22_X2 U8906 ( .A1(n26389), .A2(n26894), .B1(n25811), .B2(n15930), .ZN(
        n24123) );
  OAI22_X2 U8908 ( .A1(n26389), .A2(n26895), .B1(n25808), .B2(n15930), .ZN(
        n24124) );
  OAI22_X2 U8910 ( .A1(n26389), .A2(n26896), .B1(n25805), .B2(n15930), .ZN(
        n24125) );
  OAI22_X2 U8912 ( .A1(n26389), .A2(n26897), .B1(n25802), .B2(n15930), .ZN(
        n24126) );
  OAI22_X2 U8914 ( .A1(n26389), .A2(n26898), .B1(n25798), .B2(n15930), .ZN(
        n24127) );
  OAI22_X2 U8916 ( .A1(n26389), .A2(n26899), .B1(n25793), .B2(n15930), .ZN(
        n24128) );
  OAI22_X2 U8918 ( .A1(n26389), .A2(n26900), .B1(n25790), .B2(n15930), .ZN(
        n24129) );
  OAI22_X2 U8920 ( .A1(n26389), .A2(n26901), .B1(n25787), .B2(n15930), .ZN(
        n24130) );
  OAI22_X2 U8922 ( .A1(n26389), .A2(n26902), .B1(n25784), .B2(n15930), .ZN(
        n24131) );
  OAI22_X2 U8926 ( .A1(n26388), .A2(n27143), .B1(n25833), .B2(n15947), .ZN(
        n24132) );
  OAI22_X2 U8928 ( .A1(n26388), .A2(n27144), .B1(n25829), .B2(n15947), .ZN(
        n24133) );
  OAI22_X2 U8930 ( .A1(n26388), .A2(n27145), .B1(n25825), .B2(n15947), .ZN(
        n24134) );
  OAI22_X2 U8932 ( .A1(n26388), .A2(n27146), .B1(n25822), .B2(n15947), .ZN(
        n24135) );
  OAI22_X2 U8934 ( .A1(n26388), .A2(n27147), .B1(n25819), .B2(n15947), .ZN(
        n24136) );
  OAI22_X2 U8936 ( .A1(n26388), .A2(n27148), .B1(n25816), .B2(n15947), .ZN(
        n24137) );
  OAI22_X2 U8938 ( .A1(n26388), .A2(n27149), .B1(n25813), .B2(n15947), .ZN(
        n24138) );
  OAI22_X2 U8940 ( .A1(n26388), .A2(n27150), .B1(n25810), .B2(n15947), .ZN(
        n24139) );
  OAI22_X2 U8942 ( .A1(n26388), .A2(n27151), .B1(n25807), .B2(n15947), .ZN(
        n24140) );
  OAI22_X2 U8944 ( .A1(n26388), .A2(n27152), .B1(n25804), .B2(n15947), .ZN(
        n24141) );
  OAI22_X2 U8946 ( .A1(n26388), .A2(n27153), .B1(n25801), .B2(n15947), .ZN(
        n24142) );
  OAI22_X2 U8948 ( .A1(n26388), .A2(n27154), .B1(n25798), .B2(n15947), .ZN(
        n24143) );
  OAI22_X2 U8950 ( .A1(n26388), .A2(n27155), .B1(n25793), .B2(n15947), .ZN(
        n24144) );
  OAI22_X2 U8952 ( .A1(n26388), .A2(n27156), .B1(n25789), .B2(n15947), .ZN(
        n24145) );
  OAI22_X2 U8954 ( .A1(n26388), .A2(n27157), .B1(n25786), .B2(n15947), .ZN(
        n24146) );
  OAI22_X2 U8956 ( .A1(n26388), .A2(n27158), .B1(n25783), .B2(n15947), .ZN(
        n24147) );
  OAI22_X2 U8960 ( .A1(n26387), .A2(n27399), .B1(n25832), .B2(n15949), .ZN(
        n24148) );
  OAI22_X2 U8962 ( .A1(n26387), .A2(n27400), .B1(n25829), .B2(n15949), .ZN(
        n24149) );
  OAI22_X2 U8964 ( .A1(n26387), .A2(n27401), .B1(n25824), .B2(n15949), .ZN(
        n24150) );
  OAI22_X2 U8966 ( .A1(n26387), .A2(n27402), .B1(n25821), .B2(n15949), .ZN(
        n24151) );
  OAI22_X2 U8968 ( .A1(n26387), .A2(n27403), .B1(n25818), .B2(n15949), .ZN(
        n24152) );
  OAI22_X2 U8970 ( .A1(n26387), .A2(n27404), .B1(n25815), .B2(n15949), .ZN(
        n24153) );
  OAI22_X2 U8972 ( .A1(n26387), .A2(n27405), .B1(n25812), .B2(n15949), .ZN(
        n24154) );
  OAI22_X2 U8974 ( .A1(n26387), .A2(n27406), .B1(n25809), .B2(n15949), .ZN(
        n24155) );
  OAI22_X2 U8976 ( .A1(n26387), .A2(n27407), .B1(n25806), .B2(n15949), .ZN(
        n24156) );
  OAI22_X2 U8978 ( .A1(n26387), .A2(n27408), .B1(n25803), .B2(n15949), .ZN(
        n24157) );
  OAI22_X2 U8980 ( .A1(n26387), .A2(n27409), .B1(n25800), .B2(n15949), .ZN(
        n24158) );
  OAI22_X2 U8982 ( .A1(n26387), .A2(n27410), .B1(n25798), .B2(n15949), .ZN(
        n24159) );
  OAI22_X2 U8984 ( .A1(n26387), .A2(n27411), .B1(n25793), .B2(n15949), .ZN(
        n24160) );
  OAI22_X2 U8986 ( .A1(n26387), .A2(n27412), .B1(n25788), .B2(n15949), .ZN(
        n24161) );
  OAI22_X2 U8988 ( .A1(n26387), .A2(n27413), .B1(n25785), .B2(n15949), .ZN(
        n24162) );
  OAI22_X2 U8990 ( .A1(n26387), .A2(n27414), .B1(n25782), .B2(n15949), .ZN(
        n24163) );
  NOR2_X2 U8995 ( .A1(n15950), .A2(n22381), .ZN(n15823) );
  OAI22_X2 U8996 ( .A1(n26454), .A2(n26615), .B1(n25832), .B2(n15952), .ZN(
        n24164) );
  OAI22_X2 U8998 ( .A1(n26454), .A2(n26616), .B1(n25830), .B2(n15952), .ZN(
        n24165) );
  OAI22_X2 U9000 ( .A1(n26454), .A2(n26617), .B1(n25824), .B2(n15952), .ZN(
        n24166) );
  OAI22_X2 U9002 ( .A1(n26454), .A2(n26618), .B1(n25821), .B2(n15952), .ZN(
        n24167) );
  OAI22_X2 U9004 ( .A1(n26454), .A2(n26619), .B1(n25818), .B2(n15952), .ZN(
        n24168) );
  OAI22_X2 U9006 ( .A1(n26454), .A2(n26620), .B1(n25815), .B2(n15952), .ZN(
        n24169) );
  OAI22_X2 U9008 ( .A1(n26454), .A2(n26621), .B1(n25812), .B2(n15952), .ZN(
        n24170) );
  OAI22_X2 U9010 ( .A1(n26454), .A2(n26622), .B1(n25809), .B2(n15952), .ZN(
        n24171) );
  OAI22_X2 U9012 ( .A1(n26454), .A2(n26623), .B1(n25806), .B2(n15952), .ZN(
        n24172) );
  OAI22_X2 U9014 ( .A1(n26454), .A2(n26624), .B1(n25803), .B2(n15952), .ZN(
        n24173) );
  OAI22_X2 U9016 ( .A1(n26454), .A2(n26625), .B1(n25800), .B2(n15952), .ZN(
        n24174) );
  OAI22_X2 U9018 ( .A1(n26454), .A2(n26626), .B1(n25799), .B2(n15952), .ZN(
        n24175) );
  OAI22_X2 U9020 ( .A1(n26454), .A2(n26627), .B1(n25794), .B2(n15952), .ZN(
        n24176) );
  OAI22_X2 U9022 ( .A1(n26454), .A2(n26628), .B1(n25788), .B2(n15952), .ZN(
        n24177) );
  OAI22_X2 U9024 ( .A1(n26454), .A2(n26629), .B1(n25785), .B2(n15952), .ZN(
        n24178) );
  OAI22_X2 U9026 ( .A1(n26454), .A2(n26630), .B1(n25782), .B2(n15952), .ZN(
        n24179) );
  OAI22_X2 U9030 ( .A1(n26453), .A2(n27671), .B1(n25832), .B2(n15955), .ZN(
        n24180) );
  OAI22_X2 U9032 ( .A1(n26453), .A2(n27672), .B1(n25830), .B2(n15955), .ZN(
        n24181) );
  OAI22_X2 U9034 ( .A1(n26453), .A2(n27673), .B1(n25824), .B2(n15955), .ZN(
        n24182) );
  OAI22_X2 U9036 ( .A1(n26453), .A2(n27674), .B1(n25821), .B2(n15955), .ZN(
        n24183) );
  OAI22_X2 U9038 ( .A1(n26453), .A2(n27675), .B1(n25818), .B2(n15955), .ZN(
        n24184) );
  OAI22_X2 U9040 ( .A1(n26453), .A2(n27676), .B1(n25815), .B2(n15955), .ZN(
        n24185) );
  OAI22_X2 U9042 ( .A1(n26453), .A2(n27677), .B1(n25812), .B2(n15955), .ZN(
        n24186) );
  OAI22_X2 U9044 ( .A1(n26453), .A2(n27678), .B1(n25809), .B2(n15955), .ZN(
        n24187) );
  OAI22_X2 U9046 ( .A1(n26453), .A2(n27679), .B1(n25806), .B2(n15955), .ZN(
        n24188) );
  OAI22_X2 U9048 ( .A1(n26453), .A2(n27680), .B1(n25803), .B2(n15955), .ZN(
        n24189) );
  OAI22_X2 U9050 ( .A1(n26453), .A2(n27681), .B1(n25800), .B2(n15955), .ZN(
        n24190) );
  OAI22_X2 U9052 ( .A1(n26453), .A2(n27682), .B1(n25799), .B2(n15955), .ZN(
        n24191) );
  OAI22_X2 U9054 ( .A1(n26453), .A2(n27683), .B1(n25794), .B2(n15955), .ZN(
        n24192) );
  OAI22_X2 U9056 ( .A1(n26453), .A2(n27684), .B1(n25788), .B2(n15955), .ZN(
        n24193) );
  OAI22_X2 U9058 ( .A1(n26453), .A2(n27685), .B1(n25785), .B2(n15955), .ZN(
        n24194) );
  OAI22_X2 U9060 ( .A1(n26453), .A2(n27686), .B1(n25782), .B2(n15955), .ZN(
        n24195) );
  OAI22_X2 U9064 ( .A1(n26452), .A2(n26903), .B1(n25834), .B2(n15972), .ZN(
        n24196) );
  OAI22_X2 U9066 ( .A1(n26452), .A2(n26904), .B1(n25830), .B2(n15972), .ZN(
        n24197) );
  OAI22_X2 U9068 ( .A1(n26452), .A2(n26905), .B1(n25826), .B2(n15972), .ZN(
        n24198) );
  OAI22_X2 U9070 ( .A1(n26452), .A2(n26906), .B1(n25823), .B2(n15972), .ZN(
        n24199) );
  OAI22_X2 U9072 ( .A1(n26452), .A2(n26907), .B1(n25820), .B2(n15972), .ZN(
        n24200) );
  OAI22_X2 U9074 ( .A1(n26452), .A2(n26908), .B1(n25817), .B2(n15972), .ZN(
        n24201) );
  OAI22_X2 U9076 ( .A1(n26452), .A2(n26909), .B1(n25814), .B2(n15972), .ZN(
        n24202) );
  OAI22_X2 U9078 ( .A1(n26452), .A2(n26910), .B1(n25811), .B2(n15972), .ZN(
        n24203) );
  OAI22_X2 U9080 ( .A1(n26452), .A2(n26911), .B1(n25808), .B2(n15972), .ZN(
        n24204) );
  OAI22_X2 U9082 ( .A1(n26452), .A2(n26912), .B1(n25805), .B2(n15972), .ZN(
        n24205) );
  OAI22_X2 U9084 ( .A1(n26452), .A2(n26913), .B1(n25802), .B2(n15972), .ZN(
        n24206) );
  OAI22_X2 U9086 ( .A1(n26452), .A2(n26914), .B1(n25799), .B2(n15972), .ZN(
        n24207) );
  OAI22_X2 U9088 ( .A1(n26452), .A2(n26915), .B1(n25794), .B2(n15972), .ZN(
        n24208) );
  OAI22_X2 U9090 ( .A1(n26452), .A2(n26916), .B1(n25790), .B2(n15972), .ZN(
        n24209) );
  OAI22_X2 U9092 ( .A1(n26452), .A2(n26917), .B1(n25787), .B2(n15972), .ZN(
        n24210) );
  OAI22_X2 U9094 ( .A1(n26452), .A2(n26918), .B1(n25784), .B2(n15972), .ZN(
        n24211) );
  OAI22_X2 U9098 ( .A1(n26451), .A2(n27159), .B1(n25833), .B2(n15974), .ZN(
        n24212) );
  OAI22_X2 U9100 ( .A1(n26451), .A2(n27160), .B1(n25830), .B2(n15974), .ZN(
        n24213) );
  OAI22_X2 U9102 ( .A1(n26451), .A2(n27161), .B1(n25825), .B2(n15974), .ZN(
        n24214) );
  OAI22_X2 U9104 ( .A1(n26451), .A2(n27162), .B1(n25822), .B2(n15974), .ZN(
        n24215) );
  OAI22_X2 U9106 ( .A1(n26451), .A2(n27163), .B1(n25819), .B2(n15974), .ZN(
        n24216) );
  OAI22_X2 U9108 ( .A1(n26451), .A2(n27164), .B1(n25816), .B2(n15974), .ZN(
        n24217) );
  OAI22_X2 U9110 ( .A1(n26451), .A2(n27165), .B1(n25813), .B2(n15974), .ZN(
        n24218) );
  OAI22_X2 U9112 ( .A1(n26451), .A2(n27166), .B1(n25810), .B2(n15974), .ZN(
        n24219) );
  OAI22_X2 U9114 ( .A1(n26451), .A2(n27167), .B1(n25807), .B2(n15974), .ZN(
        n24220) );
  OAI22_X2 U9116 ( .A1(n26451), .A2(n27168), .B1(n25804), .B2(n15974), .ZN(
        n24221) );
  OAI22_X2 U9118 ( .A1(n26451), .A2(n27169), .B1(n25801), .B2(n15974), .ZN(
        n24222) );
  OAI22_X2 U9120 ( .A1(n26451), .A2(n27170), .B1(n25799), .B2(n15974), .ZN(
        n24223) );
  OAI22_X2 U9122 ( .A1(n26451), .A2(n27171), .B1(n25794), .B2(n15974), .ZN(
        n24224) );
  OAI22_X2 U9124 ( .A1(n26451), .A2(n27172), .B1(n25789), .B2(n15974), .ZN(
        n24225) );
  OAI22_X2 U9126 ( .A1(n26451), .A2(n27173), .B1(n25786), .B2(n15974), .ZN(
        n24226) );
  OAI22_X2 U9128 ( .A1(n26451), .A2(n27174), .B1(n25783), .B2(n15974), .ZN(
        n24227) );
  OAI22_X2 U9132 ( .A1(n26450), .A2(n27415), .B1(n25832), .B2(n15976), .ZN(
        n24228) );
  OAI22_X2 U9134 ( .A1(n26450), .A2(n27416), .B1(n25830), .B2(n15976), .ZN(
        n24229) );
  OAI22_X2 U9136 ( .A1(n26450), .A2(n27417), .B1(n25824), .B2(n15976), .ZN(
        n24230) );
  OAI22_X2 U9138 ( .A1(n26450), .A2(n27418), .B1(n25821), .B2(n15976), .ZN(
        n24231) );
  OAI22_X2 U9140 ( .A1(n26450), .A2(n27419), .B1(n25818), .B2(n15976), .ZN(
        n24232) );
  OAI22_X2 U9142 ( .A1(n26450), .A2(n27420), .B1(n25815), .B2(n15976), .ZN(
        n24233) );
  OAI22_X2 U9144 ( .A1(n26450), .A2(n27421), .B1(n25812), .B2(n15976), .ZN(
        n24234) );
  OAI22_X2 U9146 ( .A1(n26450), .A2(n27422), .B1(n25809), .B2(n15976), .ZN(
        n24235) );
  OAI22_X2 U9148 ( .A1(n26450), .A2(n27423), .B1(n25806), .B2(n15976), .ZN(
        n24236) );
  OAI22_X2 U9150 ( .A1(n26450), .A2(n27424), .B1(n25803), .B2(n15976), .ZN(
        n24237) );
  OAI22_X2 U9152 ( .A1(n26450), .A2(n27425), .B1(n25800), .B2(n15976), .ZN(
        n24238) );
  OAI22_X2 U9154 ( .A1(n26450), .A2(n27426), .B1(n25799), .B2(n15976), .ZN(
        n24239) );
  OAI22_X2 U9156 ( .A1(n26450), .A2(n27427), .B1(n25794), .B2(n15976), .ZN(
        n24240) );
  OAI22_X2 U9158 ( .A1(n26450), .A2(n27428), .B1(n25788), .B2(n15976), .ZN(
        n24241) );
  OAI22_X2 U9160 ( .A1(n26450), .A2(n27429), .B1(n25785), .B2(n15976), .ZN(
        n24242) );
  OAI22_X2 U9162 ( .A1(n26450), .A2(n27430), .B1(n25782), .B2(n15976), .ZN(
        n24243) );
  OAI22_X2 U9167 ( .A1(n26445), .A2(n26743), .B1(n25834), .B2(n15979), .ZN(
        n24244) );
  OAI22_X2 U9169 ( .A1(n26445), .A2(n26744), .B1(n25830), .B2(n15979), .ZN(
        n24245) );
  OAI22_X2 U9171 ( .A1(n26445), .A2(n26745), .B1(n25826), .B2(n15979), .ZN(
        n24246) );
  OAI22_X2 U9173 ( .A1(n26445), .A2(n26746), .B1(n25823), .B2(n15979), .ZN(
        n24247) );
  OAI22_X2 U9175 ( .A1(n26445), .A2(n26747), .B1(n25820), .B2(n15979), .ZN(
        n24248) );
  OAI22_X2 U9177 ( .A1(n26445), .A2(n26748), .B1(n25817), .B2(n15979), .ZN(
        n24249) );
  OAI22_X2 U9179 ( .A1(n26445), .A2(n26749), .B1(n25814), .B2(n15979), .ZN(
        n24250) );
  OAI22_X2 U9181 ( .A1(n26445), .A2(n26750), .B1(n25811), .B2(n15979), .ZN(
        n24251) );
  OAI22_X2 U9183 ( .A1(n26445), .A2(n26751), .B1(n25808), .B2(n15979), .ZN(
        n24252) );
  OAI22_X2 U9185 ( .A1(n26445), .A2(n26752), .B1(n25805), .B2(n15979), .ZN(
        n24253) );
  OAI22_X2 U9187 ( .A1(n26445), .A2(n26753), .B1(n25802), .B2(n15979), .ZN(
        n24254) );
  OAI22_X2 U9189 ( .A1(n26445), .A2(n26754), .B1(n25799), .B2(n15979), .ZN(
        n24255) );
  OAI22_X2 U9191 ( .A1(n26445), .A2(n26755), .B1(n25794), .B2(n15979), .ZN(
        n24256) );
  OAI22_X2 U9193 ( .A1(n26445), .A2(n26756), .B1(n25790), .B2(n15979), .ZN(
        n24257) );
  OAI22_X2 U9195 ( .A1(n26445), .A2(n26757), .B1(n25787), .B2(n15979), .ZN(
        n24258) );
  OAI22_X2 U9197 ( .A1(n26445), .A2(n26758), .B1(n25784), .B2(n15979), .ZN(
        n24259) );
  OAI22_X2 U9201 ( .A1(n26444), .A2(n27687), .B1(n25834), .B2(n15982), .ZN(
        n24260) );
  OAI22_X2 U9203 ( .A1(n26444), .A2(n27688), .B1(n25830), .B2(n15982), .ZN(
        n24261) );
  OAI22_X2 U9205 ( .A1(n26444), .A2(n27689), .B1(n25826), .B2(n15982), .ZN(
        n24262) );
  OAI22_X2 U9207 ( .A1(n26444), .A2(n27690), .B1(n25823), .B2(n15982), .ZN(
        n24263) );
  OAI22_X2 U9209 ( .A1(n26444), .A2(n27691), .B1(n25820), .B2(n15982), .ZN(
        n24264) );
  OAI22_X2 U9211 ( .A1(n26444), .A2(n27692), .B1(n25817), .B2(n15982), .ZN(
        n24265) );
  OAI22_X2 U9213 ( .A1(n26444), .A2(n27693), .B1(n25814), .B2(n15982), .ZN(
        n24266) );
  OAI22_X2 U9215 ( .A1(n26444), .A2(n27694), .B1(n25811), .B2(n15982), .ZN(
        n24267) );
  OAI22_X2 U9217 ( .A1(n26444), .A2(n27695), .B1(n25808), .B2(n15982), .ZN(
        n24268) );
  OAI22_X2 U9219 ( .A1(n26444), .A2(n27696), .B1(n25805), .B2(n15982), .ZN(
        n24269) );
  OAI22_X2 U9221 ( .A1(n26444), .A2(n27697), .B1(n25802), .B2(n15982), .ZN(
        n24270) );
  OAI22_X2 U9223 ( .A1(n26444), .A2(n27698), .B1(n25799), .B2(n15982), .ZN(
        n24271) );
  OAI22_X2 U9225 ( .A1(n26444), .A2(n27699), .B1(n25794), .B2(n15982), .ZN(
        n24272) );
  OAI22_X2 U9227 ( .A1(n26444), .A2(n27700), .B1(n25790), .B2(n15982), .ZN(
        n24273) );
  OAI22_X2 U9229 ( .A1(n26444), .A2(n27701), .B1(n25787), .B2(n15982), .ZN(
        n24274) );
  OAI22_X2 U9231 ( .A1(n26444), .A2(n27702), .B1(n25784), .B2(n15982), .ZN(
        n24275) );
  OAI22_X2 U9235 ( .A1(n26443), .A2(n26919), .B1(n25833), .B2(n15999), .ZN(
        n24276) );
  OAI22_X2 U9237 ( .A1(n26443), .A2(n26920), .B1(n25830), .B2(n15999), .ZN(
        n24277) );
  OAI22_X2 U9239 ( .A1(n26443), .A2(n26921), .B1(n25825), .B2(n15999), .ZN(
        n24278) );
  OAI22_X2 U9241 ( .A1(n26443), .A2(n26922), .B1(n25822), .B2(n15999), .ZN(
        n24279) );
  OAI22_X2 U9243 ( .A1(n26443), .A2(n26923), .B1(n25819), .B2(n15999), .ZN(
        n24280) );
  OAI22_X2 U9245 ( .A1(n26443), .A2(n26924), .B1(n25816), .B2(n15999), .ZN(
        n24281) );
  OAI22_X2 U9247 ( .A1(n26443), .A2(n26925), .B1(n25813), .B2(n15999), .ZN(
        n24282) );
  OAI22_X2 U9249 ( .A1(n26443), .A2(n26926), .B1(n25810), .B2(n15999), .ZN(
        n24283) );
  OAI22_X2 U9251 ( .A1(n26443), .A2(n26927), .B1(n25807), .B2(n15999), .ZN(
        n24284) );
  OAI22_X2 U9253 ( .A1(n26443), .A2(n26928), .B1(n25804), .B2(n15999), .ZN(
        n24285) );
  OAI22_X2 U9255 ( .A1(n26443), .A2(n26929), .B1(n25801), .B2(n15999), .ZN(
        n24286) );
  OAI22_X2 U9257 ( .A1(n26443), .A2(n26930), .B1(n25799), .B2(n15999), .ZN(
        n24287) );
  OAI22_X2 U9259 ( .A1(n26443), .A2(n26931), .B1(n25794), .B2(n15999), .ZN(
        n24288) );
  OAI22_X2 U9261 ( .A1(n26443), .A2(n26932), .B1(n25789), .B2(n15999), .ZN(
        n24289) );
  OAI22_X2 U9263 ( .A1(n26443), .A2(n26933), .B1(n25786), .B2(n15999), .ZN(
        n24290) );
  OAI22_X2 U9265 ( .A1(n26443), .A2(n26934), .B1(n25783), .B2(n15999), .ZN(
        n24291) );
  OAI22_X2 U9269 ( .A1(n26442), .A2(n27175), .B1(n25832), .B2(n16001), .ZN(
        n24292) );
  OAI22_X2 U9271 ( .A1(n26442), .A2(n27176), .B1(n25830), .B2(n16001), .ZN(
        n24293) );
  OAI22_X2 U9273 ( .A1(n26442), .A2(n27177), .B1(n25824), .B2(n16001), .ZN(
        n24294) );
  OAI22_X2 U9275 ( .A1(n26442), .A2(n27178), .B1(n25821), .B2(n16001), .ZN(
        n24295) );
  OAI22_X2 U9277 ( .A1(n26442), .A2(n27179), .B1(n25818), .B2(n16001), .ZN(
        n24296) );
  OAI22_X2 U9279 ( .A1(n26442), .A2(n27180), .B1(n25815), .B2(n16001), .ZN(
        n24297) );
  OAI22_X2 U9281 ( .A1(n26442), .A2(n27181), .B1(n25812), .B2(n16001), .ZN(
        n24298) );
  OAI22_X2 U9283 ( .A1(n26442), .A2(n27182), .B1(n25809), .B2(n16001), .ZN(
        n24299) );
  OAI22_X2 U9285 ( .A1(n26442), .A2(n27183), .B1(n25806), .B2(n16001), .ZN(
        n24300) );
  OAI22_X2 U9287 ( .A1(n26442), .A2(n27184), .B1(n25803), .B2(n16001), .ZN(
        n24301) );
  OAI22_X2 U9289 ( .A1(n26442), .A2(n27185), .B1(n25800), .B2(n16001), .ZN(
        n24302) );
  OAI22_X2 U9291 ( .A1(n26442), .A2(n27186), .B1(n25799), .B2(n16001), .ZN(
        n24303) );
  OAI22_X2 U9293 ( .A1(n26442), .A2(n27187), .B1(n25794), .B2(n16001), .ZN(
        n24304) );
  OAI22_X2 U9295 ( .A1(n26442), .A2(n27188), .B1(n25788), .B2(n16001), .ZN(
        n24305) );
  OAI22_X2 U9297 ( .A1(n26442), .A2(n27189), .B1(n25785), .B2(n16001), .ZN(
        n24306) );
  OAI22_X2 U9299 ( .A1(n26442), .A2(n27190), .B1(n25782), .B2(n16001), .ZN(
        n24307) );
  OAI22_X2 U9303 ( .A1(n26441), .A2(n27431), .B1(n25834), .B2(n16003), .ZN(
        n24308) );
  OAI22_X2 U9305 ( .A1(n26441), .A2(n27432), .B1(n25830), .B2(n16003), .ZN(
        n24309) );
  OAI22_X2 U9307 ( .A1(n26441), .A2(n27433), .B1(n25826), .B2(n16003), .ZN(
        n24310) );
  OAI22_X2 U9309 ( .A1(n26441), .A2(n27434), .B1(n25823), .B2(n16003), .ZN(
        n24311) );
  OAI22_X2 U9311 ( .A1(n26441), .A2(n27435), .B1(n25820), .B2(n16003), .ZN(
        n24312) );
  OAI22_X2 U9313 ( .A1(n26441), .A2(n27436), .B1(n25817), .B2(n16003), .ZN(
        n24313) );
  OAI22_X2 U9315 ( .A1(n26441), .A2(n27437), .B1(n25814), .B2(n16003), .ZN(
        n24314) );
  OAI22_X2 U9317 ( .A1(n26441), .A2(n27438), .B1(n25811), .B2(n16003), .ZN(
        n24315) );
  OAI22_X2 U9319 ( .A1(n26441), .A2(n27439), .B1(n25808), .B2(n16003), .ZN(
        n24316) );
  OAI22_X2 U9321 ( .A1(n26441), .A2(n27440), .B1(n25805), .B2(n16003), .ZN(
        n24317) );
  OAI22_X2 U9323 ( .A1(n26441), .A2(n27441), .B1(n25802), .B2(n16003), .ZN(
        n24318) );
  OAI22_X2 U9325 ( .A1(n26441), .A2(n27442), .B1(n25799), .B2(n16003), .ZN(
        n24319) );
  OAI22_X2 U9327 ( .A1(n26441), .A2(n27443), .B1(n25794), .B2(n16003), .ZN(
        n24320) );
  OAI22_X2 U9329 ( .A1(n26441), .A2(n27444), .B1(n25790), .B2(n16003), .ZN(
        n24321) );
  OAI22_X2 U9331 ( .A1(n26441), .A2(n27445), .B1(n25787), .B2(n16003), .ZN(
        n24322) );
  OAI22_X2 U9333 ( .A1(n26441), .A2(n27446), .B1(n25784), .B2(n16003), .ZN(
        n24323) );
  OAI22_X2 U9338 ( .A1(n26436), .A2(n26679), .B1(n25833), .B2(n16005), .ZN(
        n24324) );
  OAI22_X2 U9340 ( .A1(n26436), .A2(n26680), .B1(n25830), .B2(n16005), .ZN(
        n24325) );
  OAI22_X2 U9342 ( .A1(n26436), .A2(n26681), .B1(n25825), .B2(n16005), .ZN(
        n24326) );
  OAI22_X2 U9344 ( .A1(n26436), .A2(n26682), .B1(n25822), .B2(n16005), .ZN(
        n24327) );
  OAI22_X2 U9346 ( .A1(n26436), .A2(n26683), .B1(n25819), .B2(n16005), .ZN(
        n24328) );
  OAI22_X2 U9348 ( .A1(n26436), .A2(n26684), .B1(n25816), .B2(n16005), .ZN(
        n24329) );
  OAI22_X2 U9350 ( .A1(n26436), .A2(n26685), .B1(n25813), .B2(n16005), .ZN(
        n24330) );
  OAI22_X2 U9352 ( .A1(n26436), .A2(n26686), .B1(n25810), .B2(n16005), .ZN(
        n24331) );
  OAI22_X2 U9354 ( .A1(n26436), .A2(n26687), .B1(n25807), .B2(n16005), .ZN(
        n24332) );
  OAI22_X2 U9356 ( .A1(n26436), .A2(n26688), .B1(n25804), .B2(n16005), .ZN(
        n24333) );
  OAI22_X2 U9358 ( .A1(n26436), .A2(n26689), .B1(n25801), .B2(n16005), .ZN(
        n24334) );
  OAI22_X2 U9360 ( .A1(n26436), .A2(n26690), .B1(n25799), .B2(n16005), .ZN(
        n24335) );
  OAI22_X2 U9362 ( .A1(n26436), .A2(n26691), .B1(n25794), .B2(n16005), .ZN(
        n24336) );
  OAI22_X2 U9364 ( .A1(n26436), .A2(n26692), .B1(n25789), .B2(n16005), .ZN(
        n24337) );
  OAI22_X2 U9366 ( .A1(n26436), .A2(n26693), .B1(n25786), .B2(n16005), .ZN(
        n24338) );
  OAI22_X2 U9368 ( .A1(n26436), .A2(n26694), .B1(n25783), .B2(n16005), .ZN(
        n24339) );
  OAI22_X2 U9372 ( .A1(n26435), .A2(n27703), .B1(n25833), .B2(n16008), .ZN(
        n24340) );
  OAI22_X2 U9374 ( .A1(n26435), .A2(n27704), .B1(n25830), .B2(n16008), .ZN(
        n24341) );
  OAI22_X2 U9376 ( .A1(n26435), .A2(n27705), .B1(n25825), .B2(n16008), .ZN(
        n24342) );
  OAI22_X2 U9378 ( .A1(n26435), .A2(n27706), .B1(n25822), .B2(n16008), .ZN(
        n24343) );
  OAI22_X2 U9380 ( .A1(n26435), .A2(n27707), .B1(n25819), .B2(n16008), .ZN(
        n24344) );
  OAI22_X2 U9382 ( .A1(n26435), .A2(n27708), .B1(n25816), .B2(n16008), .ZN(
        n24345) );
  OAI22_X2 U9384 ( .A1(n26435), .A2(n27709), .B1(n25813), .B2(n16008), .ZN(
        n24346) );
  OAI22_X2 U9386 ( .A1(n26435), .A2(n27710), .B1(n25810), .B2(n16008), .ZN(
        n24347) );
  OAI22_X2 U9388 ( .A1(n26435), .A2(n27711), .B1(n25807), .B2(n16008), .ZN(
        n24348) );
  OAI22_X2 U9390 ( .A1(n26435), .A2(n27712), .B1(n25804), .B2(n16008), .ZN(
        n24349) );
  OAI22_X2 U9392 ( .A1(n26435), .A2(n27713), .B1(n25801), .B2(n16008), .ZN(
        n24350) );
  OAI22_X2 U9394 ( .A1(n26435), .A2(n27714), .B1(n25799), .B2(n16008), .ZN(
        n24351) );
  OAI22_X2 U9396 ( .A1(n26435), .A2(n27715), .B1(n25794), .B2(n16008), .ZN(
        n24352) );
  OAI22_X2 U9398 ( .A1(n26435), .A2(n27716), .B1(n25789), .B2(n16008), .ZN(
        n24353) );
  OAI22_X2 U9400 ( .A1(n26435), .A2(n27717), .B1(n25786), .B2(n16008), .ZN(
        n24354) );
  OAI22_X2 U9402 ( .A1(n26435), .A2(n27718), .B1(n25783), .B2(n16008), .ZN(
        n24355) );
  OAI22_X2 U9406 ( .A1(n26434), .A2(n26935), .B1(n25832), .B2(n16025), .ZN(
        n24356) );
  OAI22_X2 U9408 ( .A1(n26434), .A2(n26936), .B1(n25830), .B2(n16025), .ZN(
        n24357) );
  OAI22_X2 U9410 ( .A1(n26434), .A2(n26937), .B1(n25824), .B2(n16025), .ZN(
        n24358) );
  OAI22_X2 U9412 ( .A1(n26434), .A2(n26938), .B1(n25821), .B2(n16025), .ZN(
        n24359) );
  OAI22_X2 U9414 ( .A1(n26434), .A2(n26939), .B1(n25818), .B2(n16025), .ZN(
        n24360) );
  OAI22_X2 U9416 ( .A1(n26434), .A2(n26940), .B1(n25815), .B2(n16025), .ZN(
        n24361) );
  OAI22_X2 U9418 ( .A1(n26434), .A2(n26941), .B1(n25812), .B2(n16025), .ZN(
        n24362) );
  OAI22_X2 U9420 ( .A1(n26434), .A2(n26942), .B1(n25809), .B2(n16025), .ZN(
        n24363) );
  OAI22_X2 U9422 ( .A1(n26434), .A2(n26943), .B1(n25806), .B2(n16025), .ZN(
        n24364) );
  OAI22_X2 U9424 ( .A1(n26434), .A2(n26944), .B1(n25803), .B2(n16025), .ZN(
        n24365) );
  OAI22_X2 U9426 ( .A1(n26434), .A2(n26945), .B1(n25800), .B2(n16025), .ZN(
        n24366) );
  OAI22_X2 U9428 ( .A1(n26434), .A2(n26946), .B1(n25799), .B2(n16025), .ZN(
        n24367) );
  OAI22_X2 U9430 ( .A1(n26434), .A2(n26947), .B1(n25794), .B2(n16025), .ZN(
        n24368) );
  OAI22_X2 U9432 ( .A1(n26434), .A2(n26948), .B1(n25788), .B2(n16025), .ZN(
        n24369) );
  OAI22_X2 U9434 ( .A1(n26434), .A2(n26949), .B1(n25785), .B2(n16025), .ZN(
        n24370) );
  OAI22_X2 U9436 ( .A1(n26434), .A2(n26950), .B1(n25782), .B2(n16025), .ZN(
        n24371) );
  OAI22_X2 U9440 ( .A1(n26433), .A2(n27191), .B1(n25832), .B2(n16027), .ZN(
        n24372) );
  OAI22_X2 U9442 ( .A1(n26433), .A2(n27192), .B1(n25831), .B2(n16027), .ZN(
        n24373) );
  OAI22_X2 U9444 ( .A1(n26433), .A2(n27193), .B1(n25824), .B2(n16027), .ZN(
        n24374) );
  OAI22_X2 U9446 ( .A1(n26433), .A2(n27194), .B1(n25821), .B2(n16027), .ZN(
        n24375) );
  OAI22_X2 U9448 ( .A1(n26433), .A2(n27195), .B1(n25818), .B2(n16027), .ZN(
        n24376) );
  OAI22_X2 U9450 ( .A1(n26433), .A2(n27196), .B1(n25815), .B2(n16027), .ZN(
        n24377) );
  OAI22_X2 U9452 ( .A1(n26433), .A2(n27197), .B1(n25812), .B2(n16027), .ZN(
        n24378) );
  OAI22_X2 U9454 ( .A1(n26433), .A2(n27198), .B1(n25809), .B2(n16027), .ZN(
        n24379) );
  OAI22_X2 U9456 ( .A1(n26433), .A2(n27199), .B1(n25806), .B2(n16027), .ZN(
        n24380) );
  OAI22_X2 U9458 ( .A1(n26433), .A2(n27200), .B1(n25803), .B2(n16027), .ZN(
        n24381) );
  OAI22_X2 U9460 ( .A1(n26433), .A2(n27201), .B1(n25800), .B2(n16027), .ZN(
        n24382) );
  OAI22_X2 U9462 ( .A1(n26433), .A2(n27202), .B1(n25796), .B2(n16027), .ZN(
        n24383) );
  OAI22_X2 U9464 ( .A1(n26433), .A2(n27203), .B1(n25795), .B2(n16027), .ZN(
        n24384) );
  OAI22_X2 U9466 ( .A1(n26433), .A2(n27204), .B1(n25788), .B2(n16027), .ZN(
        n24385) );
  OAI22_X2 U9468 ( .A1(n26433), .A2(n27205), .B1(n25785), .B2(n16027), .ZN(
        n24386) );
  OAI22_X2 U9470 ( .A1(n26433), .A2(n27206), .B1(n25782), .B2(n16027), .ZN(
        n24387) );
  OAI22_X2 U9474 ( .A1(n26432), .A2(n27447), .B1(n25834), .B2(n16029), .ZN(
        n24388) );
  OAI22_X2 U9476 ( .A1(n26432), .A2(n27448), .B1(n25831), .B2(n16029), .ZN(
        n24389) );
  OAI22_X2 U9478 ( .A1(n26432), .A2(n27449), .B1(n25826), .B2(n16029), .ZN(
        n24390) );
  OAI22_X2 U9480 ( .A1(n26432), .A2(n27450), .B1(n25823), .B2(n16029), .ZN(
        n24391) );
  OAI22_X2 U9482 ( .A1(n26432), .A2(n27451), .B1(n25820), .B2(n16029), .ZN(
        n24392) );
  OAI22_X2 U9484 ( .A1(n26432), .A2(n27452), .B1(n25817), .B2(n16029), .ZN(
        n24393) );
  OAI22_X2 U9486 ( .A1(n26432), .A2(n27453), .B1(n25814), .B2(n16029), .ZN(
        n24394) );
  OAI22_X2 U9488 ( .A1(n26432), .A2(n27454), .B1(n25811), .B2(n16029), .ZN(
        n24395) );
  OAI22_X2 U9490 ( .A1(n26432), .A2(n27455), .B1(n25808), .B2(n16029), .ZN(
        n24396) );
  OAI22_X2 U9492 ( .A1(n26432), .A2(n27456), .B1(n25805), .B2(n16029), .ZN(
        n24397) );
  OAI22_X2 U9494 ( .A1(n26432), .A2(n27457), .B1(n25802), .B2(n16029), .ZN(
        n24398) );
  OAI22_X2 U9496 ( .A1(n26432), .A2(n27458), .B1(n25798), .B2(n16029), .ZN(
        n24399) );
  OAI22_X2 U9498 ( .A1(n26432), .A2(n27459), .B1(n25795), .B2(n16029), .ZN(
        n24400) );
  OAI22_X2 U9500 ( .A1(n26432), .A2(n27460), .B1(n25790), .B2(n16029), .ZN(
        n24401) );
  OAI22_X2 U9502 ( .A1(n26432), .A2(n27461), .B1(n25787), .B2(n16029), .ZN(
        n24402) );
  OAI22_X2 U9504 ( .A1(n26432), .A2(n27462), .B1(n25784), .B2(n16029), .ZN(
        n24403) );
  OAI22_X2 U9509 ( .A1(n26427), .A2(n26631), .B1(n25833), .B2(n16031), .ZN(
        n24404) );
  OAI22_X2 U9511 ( .A1(n26427), .A2(n26632), .B1(n25831), .B2(n16031), .ZN(
        n24405) );
  OAI22_X2 U9513 ( .A1(n26427), .A2(n26633), .B1(n25825), .B2(n16031), .ZN(
        n24406) );
  OAI22_X2 U9515 ( .A1(n26427), .A2(n26634), .B1(n25822), .B2(n16031), .ZN(
        n24407) );
  OAI22_X2 U9517 ( .A1(n26427), .A2(n26635), .B1(n25819), .B2(n16031), .ZN(
        n24408) );
  OAI22_X2 U9519 ( .A1(n26427), .A2(n26636), .B1(n25816), .B2(n16031), .ZN(
        n24409) );
  OAI22_X2 U9521 ( .A1(n26427), .A2(n26637), .B1(n25813), .B2(n16031), .ZN(
        n24410) );
  OAI22_X2 U9523 ( .A1(n26427), .A2(n26638), .B1(n25810), .B2(n16031), .ZN(
        n24411) );
  OAI22_X2 U9525 ( .A1(n26427), .A2(n26639), .B1(n25807), .B2(n16031), .ZN(
        n24412) );
  OAI22_X2 U9527 ( .A1(n26427), .A2(n26640), .B1(n25804), .B2(n16031), .ZN(
        n24413) );
  OAI22_X2 U9529 ( .A1(n26427), .A2(n26641), .B1(n25801), .B2(n16031), .ZN(
        n24414) );
  OAI22_X2 U9531 ( .A1(n26427), .A2(n26642), .B1(n25799), .B2(n16031), .ZN(
        n24415) );
  OAI22_X2 U9533 ( .A1(n26427), .A2(n26643), .B1(n25795), .B2(n16031), .ZN(
        n24416) );
  OAI22_X2 U9535 ( .A1(n26427), .A2(n26644), .B1(n25789), .B2(n16031), .ZN(
        n24417) );
  OAI22_X2 U9537 ( .A1(n26427), .A2(n26645), .B1(n25786), .B2(n16031), .ZN(
        n24418) );
  OAI22_X2 U9539 ( .A1(n26427), .A2(n26646), .B1(n25783), .B2(n16031), .ZN(
        n24419) );
  OAI22_X2 U9543 ( .A1(n26426), .A2(n27719), .B1(n25834), .B2(n16034), .ZN(
        n24420) );
  OAI22_X2 U9545 ( .A1(n26426), .A2(n27720), .B1(n25831), .B2(n16034), .ZN(
        n24421) );
  OAI22_X2 U9547 ( .A1(n26426), .A2(n27721), .B1(n25826), .B2(n16034), .ZN(
        n24422) );
  OAI22_X2 U9549 ( .A1(n26426), .A2(n27722), .B1(n25823), .B2(n16034), .ZN(
        n24423) );
  OAI22_X2 U9551 ( .A1(n26426), .A2(n27723), .B1(n25820), .B2(n16034), .ZN(
        n24424) );
  OAI22_X2 U9553 ( .A1(n26426), .A2(n27724), .B1(n25817), .B2(n16034), .ZN(
        n24425) );
  OAI22_X2 U9555 ( .A1(n26426), .A2(n27725), .B1(n25814), .B2(n16034), .ZN(
        n24426) );
  OAI22_X2 U9557 ( .A1(n26426), .A2(n27726), .B1(n25811), .B2(n16034), .ZN(
        n24427) );
  OAI22_X2 U9559 ( .A1(n26426), .A2(n27727), .B1(n25808), .B2(n16034), .ZN(
        n24428) );
  OAI22_X2 U9561 ( .A1(n26426), .A2(n27728), .B1(n25805), .B2(n16034), .ZN(
        n24429) );
  OAI22_X2 U9563 ( .A1(n26426), .A2(n27729), .B1(n25802), .B2(n16034), .ZN(
        n24430) );
  OAI22_X2 U9565 ( .A1(n26426), .A2(n27730), .B1(n25797), .B2(n16034), .ZN(
        n24431) );
  OAI22_X2 U9567 ( .A1(n26426), .A2(n27731), .B1(n25795), .B2(n16034), .ZN(
        n24432) );
  OAI22_X2 U9569 ( .A1(n26426), .A2(n27732), .B1(n25790), .B2(n16034), .ZN(
        n24433) );
  OAI22_X2 U9571 ( .A1(n26426), .A2(n27733), .B1(n25787), .B2(n16034), .ZN(
        n24434) );
  OAI22_X2 U9573 ( .A1(n26426), .A2(n27734), .B1(n25784), .B2(n16034), .ZN(
        n24435) );
  OAI22_X2 U9577 ( .A1(n26425), .A2(n26951), .B1(n25832), .B2(n16051), .ZN(
        n24436) );
  OAI22_X2 U9579 ( .A1(n26425), .A2(n26952), .B1(n25831), .B2(n16051), .ZN(
        n24437) );
  OAI22_X2 U9581 ( .A1(n26425), .A2(n26953), .B1(n25824), .B2(n16051), .ZN(
        n24438) );
  OAI22_X2 U9583 ( .A1(n26425), .A2(n26954), .B1(n25821), .B2(n16051), .ZN(
        n24439) );
  OAI22_X2 U9585 ( .A1(n26425), .A2(n26955), .B1(n25818), .B2(n16051), .ZN(
        n24440) );
  OAI22_X2 U9587 ( .A1(n26425), .A2(n26956), .B1(n25815), .B2(n16051), .ZN(
        n24441) );
  OAI22_X2 U9589 ( .A1(n26425), .A2(n26957), .B1(n25812), .B2(n16051), .ZN(
        n24442) );
  OAI22_X2 U9591 ( .A1(n26425), .A2(n26958), .B1(n25809), .B2(n16051), .ZN(
        n24443) );
  OAI22_X2 U9593 ( .A1(n26425), .A2(n26959), .B1(n25806), .B2(n16051), .ZN(
        n24444) );
  OAI22_X2 U9595 ( .A1(n26425), .A2(n26960), .B1(n25803), .B2(n16051), .ZN(
        n24445) );
  OAI22_X2 U9597 ( .A1(n26425), .A2(n26961), .B1(n25800), .B2(n16051), .ZN(
        n24446) );
  OAI22_X2 U9599 ( .A1(n26425), .A2(n26962), .B1(n25799), .B2(n16051), .ZN(
        n24447) );
  OAI22_X2 U9601 ( .A1(n26425), .A2(n26963), .B1(n25795), .B2(n16051), .ZN(
        n24448) );
  OAI22_X2 U9603 ( .A1(n26425), .A2(n26964), .B1(n25788), .B2(n16051), .ZN(
        n24449) );
  OAI22_X2 U9605 ( .A1(n26425), .A2(n26965), .B1(n25785), .B2(n16051), .ZN(
        n24450) );
  OAI22_X2 U9607 ( .A1(n26425), .A2(n26966), .B1(n25782), .B2(n16051), .ZN(
        n24451) );
  OAI22_X2 U9611 ( .A1(n26424), .A2(n27207), .B1(n25834), .B2(n16053), .ZN(
        n24452) );
  OAI22_X2 U9613 ( .A1(n26424), .A2(n27208), .B1(n25831), .B2(n16053), .ZN(
        n24453) );
  OAI22_X2 U9615 ( .A1(n26424), .A2(n27209), .B1(n25826), .B2(n16053), .ZN(
        n24454) );
  OAI22_X2 U9617 ( .A1(n26424), .A2(n27210), .B1(n25823), .B2(n16053), .ZN(
        n24455) );
  OAI22_X2 U9619 ( .A1(n26424), .A2(n27211), .B1(n25820), .B2(n16053), .ZN(
        n24456) );
  OAI22_X2 U9621 ( .A1(n26424), .A2(n27212), .B1(n25817), .B2(n16053), .ZN(
        n24457) );
  OAI22_X2 U9623 ( .A1(n26424), .A2(n27213), .B1(n25814), .B2(n16053), .ZN(
        n24458) );
  OAI22_X2 U9625 ( .A1(n26424), .A2(n27214), .B1(n25811), .B2(n16053), .ZN(
        n24459) );
  OAI22_X2 U9627 ( .A1(n26424), .A2(n27215), .B1(n25808), .B2(n16053), .ZN(
        n24460) );
  OAI22_X2 U9629 ( .A1(n26424), .A2(n27216), .B1(n25805), .B2(n16053), .ZN(
        n24461) );
  OAI22_X2 U9631 ( .A1(n26424), .A2(n27217), .B1(n25802), .B2(n16053), .ZN(
        n24462) );
  OAI22_X2 U9633 ( .A1(n26424), .A2(n27218), .B1(n25797), .B2(n16053), .ZN(
        n24463) );
  OAI22_X2 U9635 ( .A1(n26424), .A2(n27219), .B1(n25795), .B2(n16053), .ZN(
        n24464) );
  OAI22_X2 U9637 ( .A1(n26424), .A2(n27220), .B1(n25790), .B2(n16053), .ZN(
        n24465) );
  OAI22_X2 U9639 ( .A1(n26424), .A2(n27221), .B1(n25787), .B2(n16053), .ZN(
        n24466) );
  OAI22_X2 U9641 ( .A1(n26424), .A2(n27222), .B1(n25784), .B2(n16053), .ZN(
        n24467) );
  OAI22_X2 U9645 ( .A1(n26423), .A2(n27463), .B1(n25833), .B2(n16055), .ZN(
        n24468) );
  OAI22_X2 U9647 ( .A1(n26423), .A2(n27464), .B1(n25831), .B2(n16055), .ZN(
        n24469) );
  OAI22_X2 U9649 ( .A1(n26423), .A2(n27465), .B1(n25825), .B2(n16055), .ZN(
        n24470) );
  OAI22_X2 U9651 ( .A1(n26423), .A2(n27466), .B1(n25822), .B2(n16055), .ZN(
        n24471) );
  OAI22_X2 U9653 ( .A1(n26423), .A2(n27467), .B1(n25819), .B2(n16055), .ZN(
        n24472) );
  OAI22_X2 U9655 ( .A1(n26423), .A2(n27468), .B1(n25816), .B2(n16055), .ZN(
        n24473) );
  OAI22_X2 U9657 ( .A1(n26423), .A2(n27469), .B1(n25813), .B2(n16055), .ZN(
        n24474) );
  OAI22_X2 U9659 ( .A1(n26423), .A2(n27470), .B1(n25810), .B2(n16055), .ZN(
        n24475) );
  OAI22_X2 U9661 ( .A1(n26423), .A2(n27471), .B1(n25807), .B2(n16055), .ZN(
        n24476) );
  OAI22_X2 U9663 ( .A1(n26423), .A2(n27472), .B1(n25804), .B2(n16055), .ZN(
        n24477) );
  OAI22_X2 U9665 ( .A1(n26423), .A2(n27473), .B1(n25801), .B2(n16055), .ZN(
        n24478) );
  OAI22_X2 U9667 ( .A1(n26423), .A2(n27474), .B1(n25799), .B2(n16055), .ZN(
        n24479) );
  OAI22_X2 U9669 ( .A1(n26423), .A2(n27475), .B1(n25795), .B2(n16055), .ZN(
        n24480) );
  OAI22_X2 U9671 ( .A1(n26423), .A2(n27476), .B1(n25789), .B2(n16055), .ZN(
        n24481) );
  OAI22_X2 U9673 ( .A1(n26423), .A2(n27477), .B1(n25786), .B2(n16055), .ZN(
        n24482) );
  OAI22_X2 U9675 ( .A1(n26423), .A2(n27478), .B1(n25783), .B2(n16055), .ZN(
        n24483) );
  NOR2_X2 U9680 ( .A1(n26518), .A2(n22381), .ZN(n15977) );
  OAI22_X2 U9681 ( .A1(n26493), .A2(n26583), .B1(n25832), .B2(n16059), .ZN(
        n24484) );
  OAI22_X2 U9683 ( .A1(n26493), .A2(n26584), .B1(n25831), .B2(n16059), .ZN(
        n24485) );
  OAI22_X2 U9685 ( .A1(n26493), .A2(n26585), .B1(n25824), .B2(n16059), .ZN(
        n24486) );
  OAI22_X2 U9687 ( .A1(n26493), .A2(n26586), .B1(n25821), .B2(n16059), .ZN(
        n24487) );
  OAI22_X2 U9689 ( .A1(n26493), .A2(n26587), .B1(n25818), .B2(n16059), .ZN(
        n24488) );
  OAI22_X2 U9691 ( .A1(n26493), .A2(n26588), .B1(n25815), .B2(n16059), .ZN(
        n24489) );
  OAI22_X2 U9693 ( .A1(n26493), .A2(n26589), .B1(n25812), .B2(n16059), .ZN(
        n24490) );
  OAI22_X2 U9695 ( .A1(n26493), .A2(n26590), .B1(n25809), .B2(n16059), .ZN(
        n24491) );
  OAI22_X2 U9697 ( .A1(n26493), .A2(n26591), .B1(n25806), .B2(n16059), .ZN(
        n24492) );
  OAI22_X2 U9699 ( .A1(n26493), .A2(n26592), .B1(n25803), .B2(n16059), .ZN(
        n24493) );
  OAI22_X2 U9701 ( .A1(n26493), .A2(n26593), .B1(n25800), .B2(n16059), .ZN(
        n24494) );
  OAI22_X2 U9703 ( .A1(n26493), .A2(n26594), .B1(n25797), .B2(n16059), .ZN(
        n24495) );
  OAI22_X2 U9705 ( .A1(n26493), .A2(n26595), .B1(n25795), .B2(n16059), .ZN(
        n24496) );
  OAI22_X2 U9707 ( .A1(n26493), .A2(n26596), .B1(n25788), .B2(n16059), .ZN(
        n24497) );
  OAI22_X2 U9709 ( .A1(n26493), .A2(n26597), .B1(n25785), .B2(n16059), .ZN(
        n24498) );
  OAI22_X2 U9711 ( .A1(n26493), .A2(n26598), .B1(n25782), .B2(n16059), .ZN(
        n24499) );
  OAI22_X2 U9715 ( .A1(n26492), .A2(n27735), .B1(n25833), .B2(n16076), .ZN(
        n24500) );
  OAI22_X2 U9717 ( .A1(n26492), .A2(n27736), .B1(n25831), .B2(n16076), .ZN(
        n24501) );
  OAI22_X2 U9719 ( .A1(n26492), .A2(n27737), .B1(n25825), .B2(n16076), .ZN(
        n24502) );
  OAI22_X2 U9721 ( .A1(n26492), .A2(n27738), .B1(n25822), .B2(n16076), .ZN(
        n24503) );
  OAI22_X2 U9723 ( .A1(n26492), .A2(n27739), .B1(n25819), .B2(n16076), .ZN(
        n24504) );
  OAI22_X2 U9725 ( .A1(n26492), .A2(n27740), .B1(n25816), .B2(n16076), .ZN(
        n24505) );
  OAI22_X2 U9727 ( .A1(n26492), .A2(n27741), .B1(n25813), .B2(n16076), .ZN(
        n24506) );
  OAI22_X2 U9729 ( .A1(n26492), .A2(n27742), .B1(n25810), .B2(n16076), .ZN(
        n24507) );
  OAI22_X2 U9731 ( .A1(n26492), .A2(n27743), .B1(n25807), .B2(n16076), .ZN(
        n24508) );
  OAI22_X2 U9733 ( .A1(n26492), .A2(n27744), .B1(n25804), .B2(n16076), .ZN(
        n24509) );
  OAI22_X2 U9735 ( .A1(n26492), .A2(n27745), .B1(n25801), .B2(n16076), .ZN(
        n24510) );
  OAI22_X2 U9737 ( .A1(n26492), .A2(n27746), .B1(n25796), .B2(n16076), .ZN(
        n24511) );
  OAI22_X2 U9739 ( .A1(n26492), .A2(n27747), .B1(n25795), .B2(n16076), .ZN(
        n24512) );
  OAI22_X2 U9741 ( .A1(n26492), .A2(n27748), .B1(n25789), .B2(n16076), .ZN(
        n24513) );
  OAI22_X2 U9743 ( .A1(n26492), .A2(n27749), .B1(n25786), .B2(n16076), .ZN(
        n24514) );
  OAI22_X2 U9745 ( .A1(n26492), .A2(n27750), .B1(n25783), .B2(n16076), .ZN(
        n24515) );
  OAI22_X2 U9749 ( .A1(n26491), .A2(n26967), .B1(n25834), .B2(n16078), .ZN(
        n24516) );
  OAI22_X2 U9751 ( .A1(n26491), .A2(n26968), .B1(n25831), .B2(n16078), .ZN(
        n24517) );
  OAI22_X2 U9753 ( .A1(n26491), .A2(n26969), .B1(n25826), .B2(n16078), .ZN(
        n24518) );
  OAI22_X2 U9755 ( .A1(n26491), .A2(n26970), .B1(n25823), .B2(n16078), .ZN(
        n24519) );
  OAI22_X2 U9757 ( .A1(n26491), .A2(n26971), .B1(n25820), .B2(n16078), .ZN(
        n24520) );
  OAI22_X2 U9759 ( .A1(n26491), .A2(n26972), .B1(n25817), .B2(n16078), .ZN(
        n24521) );
  OAI22_X2 U9761 ( .A1(n26491), .A2(n26973), .B1(n25814), .B2(n16078), .ZN(
        n24522) );
  OAI22_X2 U9763 ( .A1(n26491), .A2(n26974), .B1(n25811), .B2(n16078), .ZN(
        n24523) );
  OAI22_X2 U9765 ( .A1(n26491), .A2(n26975), .B1(n25808), .B2(n16078), .ZN(
        n24524) );
  OAI22_X2 U9767 ( .A1(n26491), .A2(n26976), .B1(n25805), .B2(n16078), .ZN(
        n24525) );
  OAI22_X2 U9769 ( .A1(n26491), .A2(n26977), .B1(n25802), .B2(n16078), .ZN(
        n24526) );
  OAI22_X2 U9771 ( .A1(n26491), .A2(n26978), .B1(n25799), .B2(n16078), .ZN(
        n24527) );
  OAI22_X2 U9773 ( .A1(n26491), .A2(n26979), .B1(n25795), .B2(n16078), .ZN(
        n24528) );
  OAI22_X2 U9775 ( .A1(n26491), .A2(n26980), .B1(n25790), .B2(n16078), .ZN(
        n24529) );
  OAI22_X2 U9777 ( .A1(n26491), .A2(n26981), .B1(n25787), .B2(n16078), .ZN(
        n24530) );
  OAI22_X2 U9779 ( .A1(n26491), .A2(n26982), .B1(n25784), .B2(n16078), .ZN(
        n24531) );
  OAI22_X2 U9783 ( .A1(n26490), .A2(n27223), .B1(n25833), .B2(n16081), .ZN(
        n24532) );
  OAI22_X2 U9785 ( .A1(n26490), .A2(n27224), .B1(n25831), .B2(n16081), .ZN(
        n24533) );
  OAI22_X2 U9787 ( .A1(n26490), .A2(n27225), .B1(n25825), .B2(n16081), .ZN(
        n24534) );
  OAI22_X2 U9789 ( .A1(n26490), .A2(n27226), .B1(n25822), .B2(n16081), .ZN(
        n24535) );
  OAI22_X2 U9791 ( .A1(n26490), .A2(n27227), .B1(n25819), .B2(n16081), .ZN(
        n24536) );
  OAI22_X2 U9793 ( .A1(n26490), .A2(n27228), .B1(n25816), .B2(n16081), .ZN(
        n24537) );
  OAI22_X2 U9795 ( .A1(n26490), .A2(n27229), .B1(n25813), .B2(n16081), .ZN(
        n24538) );
  OAI22_X2 U9797 ( .A1(n26490), .A2(n27230), .B1(n25810), .B2(n16081), .ZN(
        n24539) );
  OAI22_X2 U9799 ( .A1(n26490), .A2(n27231), .B1(n25807), .B2(n16081), .ZN(
        n24540) );
  OAI22_X2 U9801 ( .A1(n26490), .A2(n27232), .B1(n25804), .B2(n16081), .ZN(
        n24541) );
  OAI22_X2 U9803 ( .A1(n26490), .A2(n27233), .B1(n25801), .B2(n16081), .ZN(
        n24542) );
  OAI22_X2 U9805 ( .A1(n26490), .A2(n27234), .B1(n25796), .B2(n16081), .ZN(
        n24543) );
  OAI22_X2 U9807 ( .A1(n26490), .A2(n27235), .B1(n25795), .B2(n16081), .ZN(
        n24544) );
  OAI22_X2 U9809 ( .A1(n26490), .A2(n27236), .B1(n25789), .B2(n16081), .ZN(
        n24545) );
  OAI22_X2 U9811 ( .A1(n26490), .A2(n27237), .B1(n25786), .B2(n16081), .ZN(
        n24546) );
  OAI22_X2 U9813 ( .A1(n26490), .A2(n27238), .B1(n25783), .B2(n16081), .ZN(
        n24547) );
  OAI22_X2 U9817 ( .A1(n26489), .A2(n27479), .B1(n25832), .B2(n16099), .ZN(
        n24548) );
  OAI22_X2 U9819 ( .A1(n26489), .A2(n27480), .B1(n25831), .B2(n16099), .ZN(
        n24549) );
  OAI22_X2 U9821 ( .A1(n26489), .A2(n27481), .B1(n25824), .B2(n16099), .ZN(
        n24550) );
  OAI22_X2 U9823 ( .A1(n26489), .A2(n27482), .B1(n25821), .B2(n16099), .ZN(
        n24551) );
  OAI22_X2 U9825 ( .A1(n26489), .A2(n27483), .B1(n25818), .B2(n16099), .ZN(
        n24552) );
  OAI22_X2 U9827 ( .A1(n26489), .A2(n27484), .B1(n25815), .B2(n16099), .ZN(
        n24553) );
  OAI22_X2 U9829 ( .A1(n26489), .A2(n27485), .B1(n25812), .B2(n16099), .ZN(
        n24554) );
  OAI22_X2 U9831 ( .A1(n26489), .A2(n27486), .B1(n25809), .B2(n16099), .ZN(
        n24555) );
  OAI22_X2 U9833 ( .A1(n26489), .A2(n27487), .B1(n25806), .B2(n16099), .ZN(
        n24556) );
  OAI22_X2 U9835 ( .A1(n26489), .A2(n27488), .B1(n25803), .B2(n16099), .ZN(
        n24557) );
  OAI22_X2 U9837 ( .A1(n26489), .A2(n27489), .B1(n25800), .B2(n16099), .ZN(
        n24558) );
  OAI22_X2 U9839 ( .A1(n26489), .A2(n27490), .B1(n25798), .B2(n16099), .ZN(
        n24559) );
  OAI22_X2 U9841 ( .A1(n26489), .A2(n27491), .B1(n25795), .B2(n16099), .ZN(
        n24560) );
  OAI22_X2 U9843 ( .A1(n26489), .A2(n27492), .B1(n25788), .B2(n16099), .ZN(
        n24561) );
  OAI22_X2 U9845 ( .A1(n26489), .A2(n27493), .B1(n25785), .B2(n16099), .ZN(
        n24562) );
  OAI22_X2 U9847 ( .A1(n26489), .A2(n27494), .B1(n25782), .B2(n16099), .ZN(
        n24563) );
  OAI22_X2 U9852 ( .A1(n26484), .A2(n26759), .B1(n25834), .B2(n16118), .ZN(
        n24564) );
  OAI22_X2 U9854 ( .A1(n26484), .A2(n26760), .B1(n25831), .B2(n16118), .ZN(
        n24565) );
  OAI22_X2 U9856 ( .A1(n26484), .A2(n26761), .B1(n25826), .B2(n16118), .ZN(
        n24566) );
  OAI22_X2 U9858 ( .A1(n26484), .A2(n26762), .B1(n25823), .B2(n16118), .ZN(
        n24567) );
  OAI22_X2 U9860 ( .A1(n26484), .A2(n26763), .B1(n25820), .B2(n16118), .ZN(
        n24568) );
  OAI22_X2 U9862 ( .A1(n26484), .A2(n26764), .B1(n25817), .B2(n16118), .ZN(
        n24569) );
  OAI22_X2 U9864 ( .A1(n26484), .A2(n26765), .B1(n25814), .B2(n16118), .ZN(
        n24570) );
  OAI22_X2 U9866 ( .A1(n26484), .A2(n26766), .B1(n25811), .B2(n16118), .ZN(
        n24571) );
  OAI22_X2 U9868 ( .A1(n26484), .A2(n26767), .B1(n25808), .B2(n16118), .ZN(
        n24572) );
  OAI22_X2 U9870 ( .A1(n26484), .A2(n26768), .B1(n25805), .B2(n16118), .ZN(
        n24573) );
  OAI22_X2 U9872 ( .A1(n26484), .A2(n26769), .B1(n25802), .B2(n16118), .ZN(
        n24574) );
  OAI22_X2 U9874 ( .A1(n26484), .A2(n26770), .B1(n25799), .B2(n16118), .ZN(
        n24575) );
  OAI22_X2 U9876 ( .A1(n26484), .A2(n26771), .B1(n25795), .B2(n16118), .ZN(
        n24576) );
  OAI22_X2 U9878 ( .A1(n26484), .A2(n26772), .B1(n25790), .B2(n16118), .ZN(
        n24577) );
  OAI22_X2 U9880 ( .A1(n26484), .A2(n26773), .B1(n25787), .B2(n16118), .ZN(
        n24578) );
  OAI22_X2 U9882 ( .A1(n26484), .A2(n26774), .B1(n25784), .B2(n16118), .ZN(
        n24579) );
  OAI22_X2 U9886 ( .A1(n26483), .A2(n27751), .B1(n25834), .B2(n16135), .ZN(
        n24580) );
  OAI22_X2 U9888 ( .A1(n26483), .A2(n27752), .B1(n25828), .B2(n16135), .ZN(
        n24581) );
  OAI22_X2 U9890 ( .A1(n26483), .A2(n27753), .B1(n25826), .B2(n16135), .ZN(
        n24582) );
  OAI22_X2 U9892 ( .A1(n26483), .A2(n27754), .B1(n25823), .B2(n16135), .ZN(
        n24583) );
  OAI22_X2 U9894 ( .A1(n26483), .A2(n27755), .B1(n25820), .B2(n16135), .ZN(
        n24584) );
  OAI22_X2 U9896 ( .A1(n26483), .A2(n27756), .B1(n25817), .B2(n16135), .ZN(
        n24585) );
  OAI22_X2 U9898 ( .A1(n26483), .A2(n27757), .B1(n25814), .B2(n16135), .ZN(
        n24586) );
  OAI22_X2 U9900 ( .A1(n26483), .A2(n27758), .B1(n25811), .B2(n16135), .ZN(
        n24587) );
  OAI22_X2 U9902 ( .A1(n26483), .A2(n27759), .B1(n25808), .B2(n16135), .ZN(
        n24588) );
  OAI22_X2 U9904 ( .A1(n26483), .A2(n27760), .B1(n25805), .B2(n16135), .ZN(
        n24589) );
  OAI22_X2 U9906 ( .A1(n26483), .A2(n27761), .B1(n25802), .B2(n16135), .ZN(
        n24590) );
  OAI22_X2 U9908 ( .A1(n26483), .A2(n27762), .B1(n25797), .B2(n16135), .ZN(
        n24591) );
  OAI22_X2 U9910 ( .A1(n26483), .A2(n27763), .B1(n25792), .B2(n16135), .ZN(
        n24592) );
  OAI22_X2 U9912 ( .A1(n26483), .A2(n27764), .B1(n25790), .B2(n16135), .ZN(
        n24593) );
  OAI22_X2 U9914 ( .A1(n26483), .A2(n27765), .B1(n25787), .B2(n16135), .ZN(
        n24594) );
  OAI22_X2 U9916 ( .A1(n26483), .A2(n27766), .B1(n25784), .B2(n16135), .ZN(
        n24595) );
  OAI22_X2 U9920 ( .A1(n26482), .A2(n26983), .B1(n25833), .B2(n16137), .ZN(
        n24596) );
  OAI22_X2 U9922 ( .A1(n26482), .A2(n26984), .B1(n25831), .B2(n16137), .ZN(
        n24597) );
  OAI22_X2 U9924 ( .A1(n26482), .A2(n26985), .B1(n25825), .B2(n16137), .ZN(
        n24598) );
  OAI22_X2 U9926 ( .A1(n26482), .A2(n26986), .B1(n25822), .B2(n16137), .ZN(
        n24599) );
  OAI22_X2 U9928 ( .A1(n26482), .A2(n26987), .B1(n25819), .B2(n16137), .ZN(
        n24600) );
  OAI22_X2 U9930 ( .A1(n26482), .A2(n26988), .B1(n25816), .B2(n16137), .ZN(
        n24601) );
  OAI22_X2 U9932 ( .A1(n26482), .A2(n26989), .B1(n25813), .B2(n16137), .ZN(
        n24602) );
  OAI22_X2 U9934 ( .A1(n26482), .A2(n26990), .B1(n25810), .B2(n16137), .ZN(
        n24603) );
  OAI22_X2 U9936 ( .A1(n26482), .A2(n26991), .B1(n25807), .B2(n16137), .ZN(
        n24604) );
  OAI22_X2 U9938 ( .A1(n26482), .A2(n26992), .B1(n25804), .B2(n16137), .ZN(
        n24605) );
  OAI22_X2 U9940 ( .A1(n26482), .A2(n26993), .B1(n25801), .B2(n16137), .ZN(
        n24606) );
  OAI22_X2 U9942 ( .A1(n26482), .A2(n26994), .B1(n25799), .B2(n16137), .ZN(
        n24607) );
  OAI22_X2 U9944 ( .A1(n26482), .A2(n26995), .B1(n25795), .B2(n16137), .ZN(
        n24608) );
  OAI22_X2 U9946 ( .A1(n26482), .A2(n26996), .B1(n25789), .B2(n16137), .ZN(
        n24609) );
  OAI22_X2 U9948 ( .A1(n26482), .A2(n26997), .B1(n25786), .B2(n16137), .ZN(
        n24610) );
  OAI22_X2 U9950 ( .A1(n26482), .A2(n26998), .B1(n25783), .B2(n16137), .ZN(
        n24611) );
  OAI22_X2 U9954 ( .A1(n26481), .A2(n27239), .B1(n25834), .B2(n16140), .ZN(
        n24612) );
  OAI22_X2 U9956 ( .A1(n26481), .A2(n27240), .B1(n25830), .B2(n16140), .ZN(
        n24613) );
  OAI22_X2 U9958 ( .A1(n26481), .A2(n27241), .B1(n25826), .B2(n16140), .ZN(
        n24614) );
  OAI22_X2 U9960 ( .A1(n26481), .A2(n27242), .B1(n25823), .B2(n16140), .ZN(
        n24615) );
  OAI22_X2 U9962 ( .A1(n26481), .A2(n27243), .B1(n25820), .B2(n16140), .ZN(
        n24616) );
  OAI22_X2 U9964 ( .A1(n26481), .A2(n27244), .B1(n25817), .B2(n16140), .ZN(
        n24617) );
  OAI22_X2 U9966 ( .A1(n26481), .A2(n27245), .B1(n25814), .B2(n16140), .ZN(
        n24618) );
  OAI22_X2 U9968 ( .A1(n26481), .A2(n27246), .B1(n25811), .B2(n16140), .ZN(
        n24619) );
  OAI22_X2 U9970 ( .A1(n26481), .A2(n27247), .B1(n25808), .B2(n16140), .ZN(
        n24620) );
  OAI22_X2 U9972 ( .A1(n26481), .A2(n27248), .B1(n25805), .B2(n16140), .ZN(
        n24621) );
  OAI22_X2 U9974 ( .A1(n26481), .A2(n27249), .B1(n25802), .B2(n16140), .ZN(
        n24622) );
  OAI22_X2 U9976 ( .A1(n26481), .A2(n27250), .B1(n25799), .B2(n16140), .ZN(
        n24623) );
  OAI22_X2 U9978 ( .A1(n26481), .A2(n27251), .B1(n25794), .B2(n16140), .ZN(
        n24624) );
  OAI22_X2 U9980 ( .A1(n26481), .A2(n27252), .B1(n25790), .B2(n16140), .ZN(
        n24625) );
  OAI22_X2 U9982 ( .A1(n26481), .A2(n27253), .B1(n25787), .B2(n16140), .ZN(
        n24626) );
  OAI22_X2 U9984 ( .A1(n26481), .A2(n27254), .B1(n25784), .B2(n16140), .ZN(
        n24627) );
  OAI22_X2 U9988 ( .A1(n26480), .A2(n27495), .B1(n25833), .B2(n16158), .ZN(
        n24628) );
  OAI22_X2 U9990 ( .A1(n26480), .A2(n27496), .B1(n25827), .B2(n16158), .ZN(
        n24629) );
  OAI22_X2 U9992 ( .A1(n26480), .A2(n27497), .B1(n25825), .B2(n16158), .ZN(
        n24630) );
  OAI22_X2 U9994 ( .A1(n26480), .A2(n27498), .B1(n25822), .B2(n16158), .ZN(
        n24631) );
  OAI22_X2 U9996 ( .A1(n26480), .A2(n27499), .B1(n25819), .B2(n16158), .ZN(
        n24632) );
  OAI22_X2 U9998 ( .A1(n26480), .A2(n27500), .B1(n25816), .B2(n16158), .ZN(
        n24633) );
  OAI22_X2 U10000 ( .A1(n26480), .A2(n27501), .B1(n25813), .B2(n16158), .ZN(
        n24634) );
  OAI22_X2 U10002 ( .A1(n26480), .A2(n27502), .B1(n25810), .B2(n16158), .ZN(
        n24635) );
  OAI22_X2 U10004 ( .A1(n26480), .A2(n27503), .B1(n25807), .B2(n16158), .ZN(
        n24636) );
  OAI22_X2 U10006 ( .A1(n26480), .A2(n27504), .B1(n25804), .B2(n16158), .ZN(
        n24637) );
  OAI22_X2 U10008 ( .A1(n26480), .A2(n27505), .B1(n25801), .B2(n16158), .ZN(
        n24638) );
  OAI22_X2 U10010 ( .A1(n26480), .A2(n27506), .B1(n25796), .B2(n16158), .ZN(
        n24639) );
  OAI22_X2 U10012 ( .A1(n26480), .A2(n27507), .B1(n25791), .B2(n16158), .ZN(
        n24640) );
  OAI22_X2 U10014 ( .A1(n26480), .A2(n27508), .B1(n25789), .B2(n16158), .ZN(
        n24641) );
  OAI22_X2 U10016 ( .A1(n26480), .A2(n27509), .B1(n25786), .B2(n16158), .ZN(
        n24642) );
  OAI22_X2 U10018 ( .A1(n26480), .A2(n27510), .B1(n25783), .B2(n16158), .ZN(
        n24643) );
  OAI221_X2 U10023 ( .B1(n16174), .B2(n16175), .C1(n16373), .C2(n11487), .A(
        n16176), .ZN(n24644) );
  OAI221_X2 U10025 ( .B1(n16180), .B2(n26459), .C1(n16372), .C2(n11487), .A(
        n16181), .ZN(n24645) );
  NOR2_X2 U10026 ( .A1(n11496), .A2(n16182), .ZN(n16181) );
  NOR3_X2 U10027 ( .A1(n16175), .A2(n26501), .A3(n26513), .ZN(n16182) );
  NOR3_X2 U10029 ( .A1(n12974), .A2(n16185), .A3(n16175), .ZN(n11496) );
  NAND2_X2 U10030 ( .A1(n22388), .A2(n11487), .ZN(n16175) );
  NAND2_X2 U10034 ( .A1(n26501), .A2(n16174), .ZN(n11498) );
  NAND2_X2 U10035 ( .A1(n26514), .A2(n16188), .ZN(n11497) );
  OAI22_X2 U10036 ( .A1(n16370), .A2(n11487), .B1(n12974), .B2(n16189), .ZN(
        n24646) );
  NOR2_X2 U10040 ( .A1(n13032), .A2(n26512), .ZN(n12974) );
  OAI22_X2 U10042 ( .A1(n16369), .A2(n11487), .B1(n16193), .B2(n26460), .ZN(
        n24647) );
  NAND2_X2 U10045 ( .A1(n26507), .A2(n26503), .ZN(n16194) );
  OAI221_X2 U10046 ( .B1(n16199), .B2(n26460), .C1(n16368), .C2(n11487), .A(
        n11489), .ZN(n24648) );
  NAND3_X2 U10047 ( .A1(n22387), .A2(n11487), .A3(n16200), .ZN(n11489) );
  NOR3_X2 U10050 ( .A1(n26499), .A2(n12975), .A3(n26517), .ZN(n16202) );
  NAND2_X2 U10052 ( .A1(n26503), .A2(n16196), .ZN(n11490) );
  NOR3_X2 U10053 ( .A1(n25781), .A2(n26500), .A3(n26502), .ZN(n16196) );
  NAND2_X2 U10056 ( .A1(n16188), .A2(n16192), .ZN(n11492) );
  OAI22_X2 U10057 ( .A1(n26517), .A2(n26507), .B1(n26503), .B2(n24895), .ZN(
        n16201) );
  NAND3_X2 U10060 ( .A1(n16208), .A2(n16209), .A3(n16210), .ZN(n12978) );
  OAI22_X2 U10062 ( .A1(n16366), .A2(n11487), .B1(n26460), .B2(n16211), .ZN(
        n24649) );
  NOR2_X2 U10065 ( .A1(n13032), .A2(n12889), .ZN(n12975) );
  NAND2_X2 U10066 ( .A1(n15780), .A2(n15950), .ZN(n11491) );
  NAND2_X2 U10067 ( .A1(n25252), .A2(n24895), .ZN(n15780) );
  NAND3_X2 U10068 ( .A1(n26504), .A2(n12971), .A3(n12970), .ZN(n16207) );
  NAND3_X2 U10072 ( .A1(n12972), .A2(n26504), .A3(n16210), .ZN(n16178) );
  NAND3_X2 U10074 ( .A1(n24833), .A2(n24832), .A3(n16216), .ZN(n12972) );
  NOR2_X2 U10075 ( .A1(n26505), .A2(n16177), .ZN(n16185) );
  NAND3_X2 U10076 ( .A1(n16205), .A2(n16209), .A3(n12970), .ZN(n16177) );
  NAND3_X2 U10077 ( .A1(n16218), .A2(n24832), .A3(n22386), .ZN(n12970) );
  NAND3_X2 U10078 ( .A1(n16216), .A2(n22384), .A3(n22386), .ZN(n16209) );
  NAND3_X2 U10079 ( .A1(n16218), .A2(n24833), .A3(n22384), .ZN(n16205) );
  NOR3_X2 U10081 ( .A1(n25781), .A2(n26508), .A3(n26506), .ZN(n16174) );
  OAI22_X2 U10083 ( .A1(n26475), .A2(n26695), .B1(n25832), .B2(n16221), .ZN(
        n24650) );
  OAI22_X2 U10085 ( .A1(n26475), .A2(n26696), .B1(n25828), .B2(n16221), .ZN(
        n24651) );
  OAI22_X2 U10087 ( .A1(n26475), .A2(n26697), .B1(n25824), .B2(n16221), .ZN(
        n24652) );
  OAI22_X2 U10089 ( .A1(n26475), .A2(n26698), .B1(n25821), .B2(n16221), .ZN(
        n24653) );
  OAI22_X2 U10091 ( .A1(n26475), .A2(n26699), .B1(n25818), .B2(n16221), .ZN(
        n24654) );
  OAI22_X2 U10093 ( .A1(n26475), .A2(n26700), .B1(n25815), .B2(n16221), .ZN(
        n24655) );
  OAI22_X2 U10095 ( .A1(n26475), .A2(n26701), .B1(n25812), .B2(n16221), .ZN(
        n24656) );
  OAI22_X2 U10097 ( .A1(n26475), .A2(n26702), .B1(n25809), .B2(n16221), .ZN(
        n24657) );
  OAI22_X2 U10099 ( .A1(n26475), .A2(n26703), .B1(n25806), .B2(n16221), .ZN(
        n24658) );
  OAI22_X2 U10101 ( .A1(n26475), .A2(n26704), .B1(n25803), .B2(n16221), .ZN(
        n24659) );
  OAI22_X2 U10103 ( .A1(n26475), .A2(n26705), .B1(n25800), .B2(n16221), .ZN(
        n24660) );
  OAI22_X2 U10105 ( .A1(n26475), .A2(n26706), .B1(n25797), .B2(n16221), .ZN(
        n24661) );
  OAI22_X2 U10107 ( .A1(n26475), .A2(n26707), .B1(n25792), .B2(n16221), .ZN(
        n24662) );
  OAI22_X2 U10109 ( .A1(n26475), .A2(n26708), .B1(n25788), .B2(n16221), .ZN(
        n24663) );
  OAI22_X2 U10111 ( .A1(n26475), .A2(n26709), .B1(n25785), .B2(n16221), .ZN(
        n24664) );
  OAI22_X2 U10113 ( .A1(n26475), .A2(n26710), .B1(n25782), .B2(n16221), .ZN(
        n24665) );
  OAI22_X2 U10117 ( .A1(n26474), .A2(n27767), .B1(n25832), .B2(n16238), .ZN(
        n24666) );
  OAI22_X2 U10119 ( .A1(n26474), .A2(n27768), .B1(n25831), .B2(n16238), .ZN(
        n24667) );
  OAI22_X2 U10121 ( .A1(n26474), .A2(n27769), .B1(n25824), .B2(n16238), .ZN(
        n24668) );
  OAI22_X2 U10123 ( .A1(n26474), .A2(n27770), .B1(n25821), .B2(n16238), .ZN(
        n24669) );
  OAI22_X2 U10125 ( .A1(n26474), .A2(n27771), .B1(n25818), .B2(n16238), .ZN(
        n24670) );
  OAI22_X2 U10127 ( .A1(n26474), .A2(n27772), .B1(n25815), .B2(n16238), .ZN(
        n24671) );
  OAI22_X2 U10129 ( .A1(n26474), .A2(n27773), .B1(n25812), .B2(n16238), .ZN(
        n24672) );
  OAI22_X2 U10131 ( .A1(n26474), .A2(n27774), .B1(n25809), .B2(n16238), .ZN(
        n24673) );
  OAI22_X2 U10133 ( .A1(n26474), .A2(n27775), .B1(n25806), .B2(n16238), .ZN(
        n24674) );
  OAI22_X2 U10135 ( .A1(n26474), .A2(n27776), .B1(n25803), .B2(n16238), .ZN(
        n24675) );
  OAI22_X2 U10137 ( .A1(n26474), .A2(n27777), .B1(n25800), .B2(n16238), .ZN(
        n24676) );
  OAI22_X2 U10139 ( .A1(n26474), .A2(n27778), .B1(n25797), .B2(n16238), .ZN(
        n24677) );
  OAI22_X2 U10141 ( .A1(n26474), .A2(n27779), .B1(n25795), .B2(n16238), .ZN(
        n24678) );
  OAI22_X2 U10143 ( .A1(n26474), .A2(n27780), .B1(n25788), .B2(n16238), .ZN(
        n24679) );
  OAI22_X2 U10145 ( .A1(n26474), .A2(n27781), .B1(n25785), .B2(n16238), .ZN(
        n24680) );
  OAI22_X2 U10147 ( .A1(n26474), .A2(n27782), .B1(n25782), .B2(n16238), .ZN(
        n24681) );
  OAI22_X2 U10151 ( .A1(n26473), .A2(n26999), .B1(n25834), .B2(n16240), .ZN(
        n24682) );
  OAI22_X2 U10153 ( .A1(n26473), .A2(n27000), .B1(n25830), .B2(n16240), .ZN(
        n24683) );
  OAI22_X2 U10155 ( .A1(n26473), .A2(n27001), .B1(n25826), .B2(n16240), .ZN(
        n24684) );
  OAI22_X2 U10157 ( .A1(n26473), .A2(n27002), .B1(n25823), .B2(n16240), .ZN(
        n24685) );
  OAI22_X2 U10159 ( .A1(n26473), .A2(n27003), .B1(n25820), .B2(n16240), .ZN(
        n24686) );
  OAI22_X2 U10161 ( .A1(n26473), .A2(n27004), .B1(n25817), .B2(n16240), .ZN(
        n24687) );
  OAI22_X2 U10163 ( .A1(n26473), .A2(n27005), .B1(n25814), .B2(n16240), .ZN(
        n24688) );
  OAI22_X2 U10165 ( .A1(n26473), .A2(n27006), .B1(n25811), .B2(n16240), .ZN(
        n24689) );
  OAI22_X2 U10167 ( .A1(n26473), .A2(n27007), .B1(n25808), .B2(n16240), .ZN(
        n24690) );
  OAI22_X2 U10169 ( .A1(n26473), .A2(n27008), .B1(n25805), .B2(n16240), .ZN(
        n24691) );
  OAI22_X2 U10171 ( .A1(n26473), .A2(n27009), .B1(n25802), .B2(n16240), .ZN(
        n24692) );
  OAI22_X2 U10173 ( .A1(n26473), .A2(n27010), .B1(n25799), .B2(n16240), .ZN(
        n24693) );
  OAI22_X2 U10175 ( .A1(n26473), .A2(n27011), .B1(n25794), .B2(n16240), .ZN(
        n24694) );
  OAI22_X2 U10177 ( .A1(n26473), .A2(n27012), .B1(n25790), .B2(n16240), .ZN(
        n24695) );
  OAI22_X2 U10179 ( .A1(n26473), .A2(n27013), .B1(n25787), .B2(n16240), .ZN(
        n24696) );
  OAI22_X2 U10181 ( .A1(n26473), .A2(n27014), .B1(n25784), .B2(n16240), .ZN(
        n24697) );
  OAI22_X2 U10185 ( .A1(n26472), .A2(n27255), .B1(n25832), .B2(n16243), .ZN(
        n24698) );
  OAI22_X2 U10187 ( .A1(n26472), .A2(n27256), .B1(n25827), .B2(n16243), .ZN(
        n24699) );
  OAI22_X2 U10189 ( .A1(n26472), .A2(n27257), .B1(n25824), .B2(n16243), .ZN(
        n24700) );
  OAI22_X2 U10191 ( .A1(n26472), .A2(n27258), .B1(n25821), .B2(n16243), .ZN(
        n24701) );
  OAI22_X2 U10193 ( .A1(n26472), .A2(n27259), .B1(n25818), .B2(n16243), .ZN(
        n24702) );
  OAI22_X2 U10195 ( .A1(n26472), .A2(n27260), .B1(n25815), .B2(n16243), .ZN(
        n24703) );
  OAI22_X2 U10197 ( .A1(n26472), .A2(n27261), .B1(n25812), .B2(n16243), .ZN(
        n24704) );
  OAI22_X2 U10199 ( .A1(n26472), .A2(n27262), .B1(n25809), .B2(n16243), .ZN(
        n24705) );
  OAI22_X2 U10201 ( .A1(n26472), .A2(n27263), .B1(n25806), .B2(n16243), .ZN(
        n24706) );
  OAI22_X2 U10203 ( .A1(n26472), .A2(n27264), .B1(n25803), .B2(n16243), .ZN(
        n24707) );
  OAI22_X2 U10205 ( .A1(n26472), .A2(n27265), .B1(n25800), .B2(n16243), .ZN(
        n24708) );
  OAI22_X2 U10207 ( .A1(n26472), .A2(n27266), .B1(n25796), .B2(n16243), .ZN(
        n24709) );
  OAI22_X2 U10209 ( .A1(n26472), .A2(n27267), .B1(n25791), .B2(n16243), .ZN(
        n24710) );
  OAI22_X2 U10211 ( .A1(n26472), .A2(n27268), .B1(n25788), .B2(n16243), .ZN(
        n24711) );
  OAI22_X2 U10213 ( .A1(n26472), .A2(n27269), .B1(n25785), .B2(n16243), .ZN(
        n24712) );
  OAI22_X2 U10215 ( .A1(n26472), .A2(n27270), .B1(n25782), .B2(n16243), .ZN(
        n24713) );
  OAI22_X2 U10219 ( .A1(n26471), .A2(n27511), .B1(n25834), .B2(n16261), .ZN(
        n24714) );
  OAI22_X2 U10221 ( .A1(n26471), .A2(n27512), .B1(n25828), .B2(n16261), .ZN(
        n24715) );
  OAI22_X2 U10223 ( .A1(n26471), .A2(n27513), .B1(n25826), .B2(n16261), .ZN(
        n24716) );
  OAI22_X2 U10225 ( .A1(n26471), .A2(n27514), .B1(n25823), .B2(n16261), .ZN(
        n24717) );
  OAI22_X2 U10227 ( .A1(n26471), .A2(n27515), .B1(n25820), .B2(n16261), .ZN(
        n24718) );
  OAI22_X2 U10229 ( .A1(n26471), .A2(n27516), .B1(n25817), .B2(n16261), .ZN(
        n24719) );
  OAI22_X2 U10231 ( .A1(n26471), .A2(n27517), .B1(n25814), .B2(n16261), .ZN(
        n24720) );
  OAI22_X2 U10233 ( .A1(n26471), .A2(n27518), .B1(n25811), .B2(n16261), .ZN(
        n24721) );
  OAI22_X2 U10235 ( .A1(n26471), .A2(n27519), .B1(n25808), .B2(n16261), .ZN(
        n24722) );
  OAI22_X2 U10237 ( .A1(n26471), .A2(n27520), .B1(n25805), .B2(n16261), .ZN(
        n24723) );
  OAI22_X2 U10239 ( .A1(n26471), .A2(n27521), .B1(n25802), .B2(n16261), .ZN(
        n24724) );
  OAI22_X2 U10241 ( .A1(n26471), .A2(n27522), .B1(n25797), .B2(n16261), .ZN(
        n24725) );
  OAI22_X2 U10243 ( .A1(n26471), .A2(n27523), .B1(n25792), .B2(n16261), .ZN(
        n24726) );
  OAI22_X2 U10245 ( .A1(n26471), .A2(n27524), .B1(n25790), .B2(n16261), .ZN(
        n24727) );
  OAI22_X2 U10247 ( .A1(n26471), .A2(n27525), .B1(n25787), .B2(n16261), .ZN(
        n24728) );
  OAI22_X2 U10249 ( .A1(n26471), .A2(n27526), .B1(n25784), .B2(n16261), .ZN(
        n24729) );
  NAND2_X2 U10255 ( .A1(n22389), .A2(n22390), .ZN(n16188) );
  OAI22_X2 U10256 ( .A1(n26466), .A2(n26599), .B1(n25833), .B2(n16279), .ZN(
        n24730) );
  OAI22_X2 U10258 ( .A1(n26466), .A2(n26600), .B1(n25831), .B2(n16279), .ZN(
        n24731) );
  OAI22_X2 U10260 ( .A1(n26466), .A2(n26601), .B1(n25825), .B2(n16279), .ZN(
        n24732) );
  OAI22_X2 U10262 ( .A1(n26466), .A2(n26602), .B1(n25822), .B2(n16279), .ZN(
        n24733) );
  OAI22_X2 U10264 ( .A1(n26466), .A2(n26603), .B1(n25819), .B2(n16279), .ZN(
        n24734) );
  OAI22_X2 U10266 ( .A1(n26466), .A2(n26604), .B1(n25816), .B2(n16279), .ZN(
        n24735) );
  OAI22_X2 U10268 ( .A1(n26466), .A2(n26605), .B1(n25813), .B2(n16279), .ZN(
        n24736) );
  OAI22_X2 U10270 ( .A1(n26466), .A2(n26606), .B1(n25810), .B2(n16279), .ZN(
        n24737) );
  OAI22_X2 U10272 ( .A1(n26466), .A2(n26607), .B1(n25807), .B2(n16279), .ZN(
        n24738) );
  OAI22_X2 U10274 ( .A1(n26466), .A2(n26608), .B1(n25804), .B2(n16279), .ZN(
        n24739) );
  OAI22_X2 U10276 ( .A1(n26466), .A2(n26609), .B1(n25801), .B2(n16279), .ZN(
        n24740) );
  OAI22_X2 U10278 ( .A1(n26466), .A2(n26610), .B1(n25799), .B2(n16279), .ZN(
        n24741) );
  OAI22_X2 U10280 ( .A1(n26466), .A2(n26611), .B1(n25795), .B2(n16279), .ZN(
        n24742) );
  OAI22_X2 U10282 ( .A1(n26466), .A2(n26612), .B1(n25789), .B2(n16279), .ZN(
        n24743) );
  OAI22_X2 U10284 ( .A1(n26466), .A2(n26613), .B1(n25786), .B2(n16279), .ZN(
        n24744) );
  OAI22_X2 U10286 ( .A1(n26466), .A2(n26614), .B1(n25783), .B2(n16279), .ZN(
        n24745) );
  OAI22_X2 U10290 ( .A1(n26465), .A2(n27783), .B1(n25832), .B2(n16296), .ZN(
        n24746) );
  OAI22_X2 U10292 ( .A1(n26465), .A2(n27784), .B1(n25830), .B2(n16296), .ZN(
        n24747) );
  OAI22_X2 U10294 ( .A1(n26465), .A2(n27785), .B1(n25824), .B2(n16296), .ZN(
        n24748) );
  OAI22_X2 U10296 ( .A1(n26465), .A2(n27786), .B1(n25821), .B2(n16296), .ZN(
        n24749) );
  OAI22_X2 U10298 ( .A1(n26465), .A2(n27787), .B1(n25818), .B2(n16296), .ZN(
        n24750) );
  OAI22_X2 U10300 ( .A1(n26465), .A2(n27788), .B1(n25815), .B2(n16296), .ZN(
        n24751) );
  OAI22_X2 U10302 ( .A1(n26465), .A2(n27789), .B1(n25812), .B2(n16296), .ZN(
        n24752) );
  OAI22_X2 U10304 ( .A1(n26465), .A2(n27790), .B1(n25809), .B2(n16296), .ZN(
        n24753) );
  OAI22_X2 U10306 ( .A1(n26465), .A2(n27791), .B1(n25806), .B2(n16296), .ZN(
        n24754) );
  OAI22_X2 U10308 ( .A1(n26465), .A2(n27792), .B1(n25803), .B2(n16296), .ZN(
        n24755) );
  OAI22_X2 U10310 ( .A1(n26465), .A2(n27793), .B1(n25800), .B2(n16296), .ZN(
        n24756) );
  OAI22_X2 U10312 ( .A1(n26465), .A2(n27794), .B1(n25799), .B2(n16296), .ZN(
        n24757) );
  OAI22_X2 U10314 ( .A1(n26465), .A2(n27795), .B1(n25794), .B2(n16296), .ZN(
        n24758) );
  OAI22_X2 U10316 ( .A1(n26465), .A2(n27796), .B1(n25788), .B2(n16296), .ZN(
        n24759) );
  OAI22_X2 U10318 ( .A1(n26465), .A2(n27797), .B1(n25785), .B2(n16296), .ZN(
        n24760) );
  OAI22_X2 U10320 ( .A1(n26465), .A2(n27798), .B1(n25782), .B2(n16296), .ZN(
        n24761) );
  OAI22_X2 U10325 ( .A1(n26464), .A2(n27015), .B1(n25832), .B2(n16300), .ZN(
        n24762) );
  OAI22_X2 U10327 ( .A1(n26464), .A2(n27016), .B1(n25827), .B2(n16300), .ZN(
        n24763) );
  OAI22_X2 U10329 ( .A1(n26464), .A2(n27017), .B1(n25824), .B2(n16300), .ZN(
        n24764) );
  OAI22_X2 U10331 ( .A1(n26464), .A2(n27018), .B1(n25821), .B2(n16300), .ZN(
        n24765) );
  OAI22_X2 U10333 ( .A1(n26464), .A2(n27019), .B1(n25818), .B2(n16300), .ZN(
        n24766) );
  OAI22_X2 U10335 ( .A1(n26464), .A2(n27020), .B1(n25815), .B2(n16300), .ZN(
        n24767) );
  OAI22_X2 U10337 ( .A1(n26464), .A2(n27021), .B1(n25812), .B2(n16300), .ZN(
        n24768) );
  OAI22_X2 U10339 ( .A1(n26464), .A2(n27022), .B1(n25809), .B2(n16300), .ZN(
        n24769) );
  OAI22_X2 U10341 ( .A1(n26464), .A2(n27023), .B1(n25806), .B2(n16300), .ZN(
        n24770) );
  OAI22_X2 U10343 ( .A1(n26464), .A2(n27024), .B1(n25803), .B2(n16300), .ZN(
        n24771) );
  OAI22_X2 U10345 ( .A1(n26464), .A2(n27025), .B1(n25800), .B2(n16300), .ZN(
        n24772) );
  OAI22_X2 U10347 ( .A1(n26464), .A2(n27026), .B1(n25796), .B2(n16300), .ZN(
        n24773) );
  OAI22_X2 U10349 ( .A1(n26464), .A2(n27027), .B1(n25791), .B2(n16300), .ZN(
        n24774) );
  OAI22_X2 U10351 ( .A1(n26464), .A2(n27028), .B1(n25788), .B2(n16300), .ZN(
        n24775) );
  OAI22_X2 U10353 ( .A1(n26464), .A2(n27029), .B1(n25785), .B2(n16300), .ZN(
        n24776) );
  OAI22_X2 U10355 ( .A1(n26464), .A2(n27030), .B1(n25782), .B2(n16300), .ZN(
        n24777) );
  OAI22_X2 U10360 ( .A1(n26463), .A2(n27271), .B1(n25834), .B2(n16303), .ZN(
        n24778) );
  OAI22_X2 U10362 ( .A1(n26463), .A2(n27272), .B1(n25828), .B2(n16303), .ZN(
        n24779) );
  OAI22_X2 U10364 ( .A1(n26463), .A2(n27273), .B1(n25826), .B2(n16303), .ZN(
        n24780) );
  OAI22_X2 U10366 ( .A1(n26463), .A2(n27274), .B1(n25823), .B2(n16303), .ZN(
        n24781) );
  OAI22_X2 U10368 ( .A1(n26463), .A2(n27275), .B1(n25820), .B2(n16303), .ZN(
        n24782) );
  OAI22_X2 U10370 ( .A1(n26463), .A2(n27276), .B1(n25817), .B2(n16303), .ZN(
        n24783) );
  OAI22_X2 U10372 ( .A1(n26463), .A2(n27277), .B1(n25814), .B2(n16303), .ZN(
        n24784) );
  OAI22_X2 U10374 ( .A1(n26463), .A2(n27278), .B1(n25811), .B2(n16303), .ZN(
        n24785) );
  OAI22_X2 U10376 ( .A1(n26463), .A2(n27279), .B1(n25808), .B2(n16303), .ZN(
        n24786) );
  OAI22_X2 U10378 ( .A1(n26463), .A2(n27280), .B1(n25805), .B2(n16303), .ZN(
        n24787) );
  OAI22_X2 U10380 ( .A1(n26463), .A2(n27281), .B1(n25802), .B2(n16303), .ZN(
        n24788) );
  OAI22_X2 U10382 ( .A1(n26463), .A2(n27282), .B1(n25797), .B2(n16303), .ZN(
        n24789) );
  OAI22_X2 U10384 ( .A1(n26463), .A2(n27283), .B1(n25792), .B2(n16303), .ZN(
        n24790) );
  OAI22_X2 U10386 ( .A1(n26463), .A2(n27284), .B1(n25790), .B2(n16303), .ZN(
        n24791) );
  OAI22_X2 U10388 ( .A1(n26463), .A2(n27285), .B1(n25787), .B2(n16303), .ZN(
        n24792) );
  OAI22_X2 U10390 ( .A1(n26463), .A2(n27286), .B1(n25784), .B2(n16303), .ZN(
        n24793) );
  NAND3_X2 U10395 ( .A1(n22384), .A2(n16218), .A3(n22386), .ZN(n16210) );
  OAI22_X2 U10396 ( .A1(n26462), .A2(n27527), .B1(n25833), .B2(n16321), .ZN(
        n24794) );
  OAI22_X2 U10399 ( .A1(n26462), .A2(n27528), .B1(n25830), .B2(n16321), .ZN(
        n24795) );
  OAI22_X2 U10402 ( .A1(n26462), .A2(n27529), .B1(n25825), .B2(n16321), .ZN(
        n24796) );
  OAI22_X2 U10405 ( .A1(n26462), .A2(n27530), .B1(n25822), .B2(n16321), .ZN(
        n24797) );
  OAI22_X2 U10408 ( .A1(n26462), .A2(n27531), .B1(n25819), .B2(n16321), .ZN(
        n24798) );
  OAI22_X2 U10411 ( .A1(n26462), .A2(n27532), .B1(n25816), .B2(n16321), .ZN(
        n24799) );
  OAI22_X2 U10414 ( .A1(n26462), .A2(n27533), .B1(n25813), .B2(n16321), .ZN(
        n24800) );
  OAI22_X2 U10417 ( .A1(n26462), .A2(n27534), .B1(n25810), .B2(n16321), .ZN(
        n24801) );
  OAI22_X2 U10420 ( .A1(n26462), .A2(n27535), .B1(n25807), .B2(n16321), .ZN(
        n24802) );
  OAI22_X2 U10423 ( .A1(n26462), .A2(n27536), .B1(n25804), .B2(n16321), .ZN(
        n24803) );
  OAI22_X2 U10426 ( .A1(n26462), .A2(n27537), .B1(n25801), .B2(n16321), .ZN(
        n24804) );
  OAI22_X2 U10429 ( .A1(n26462), .A2(n27538), .B1(n25799), .B2(n16321), .ZN(
        n24805) );
  OAI22_X2 U10432 ( .A1(n26462), .A2(n27539), .B1(n25794), .B2(n16321), .ZN(
        n24806) );
  OAI22_X2 U10435 ( .A1(n26462), .A2(n27540), .B1(n25789), .B2(n16321), .ZN(
        n24807) );
  OAI22_X2 U10438 ( .A1(n26462), .A2(n27541), .B1(n25786), .B2(n16321), .ZN(
        n24808) );
  OAI22_X2 U10441 ( .A1(n26462), .A2(n27542), .B1(n25783), .B2(n16321), .ZN(
        n24809) );
  NOR3_X2 U10447 ( .A1(n24895), .A2(n22381), .A3(n25252), .ZN(n16115) );
  NAND3_X2 U10450 ( .A1(n22384), .A2(n24833), .A3(n16216), .ZN(n16208) );
  NOR2_X2 U10451 ( .A1(n25400), .A2(n25249), .ZN(n16216) );
  OAI221_X2 U10452 ( .B1(n22387), .B2(n26288), .C1(n26293), .C2(n15950), .A(
        n16339), .ZN(n24810) );
  NAND3_X2 U10453 ( .A1(n16191), .A2(n13032), .A3(n26291), .ZN(n16339) );
  NOR2_X2 U10454 ( .A1(n24895), .A2(n22388), .ZN(n16191) );
  NAND2_X2 U10455 ( .A1(n22388), .A2(n24895), .ZN(n15950) );
  NAND3_X2 U10458 ( .A1(n22388), .A2(n13032), .A3(n26291), .ZN(n16341) );
  NOR2_X2 U10462 ( .A1(n22390), .A2(n22389), .ZN(n13032) );
  OAI22_X2 U10467 ( .A1(n22390), .A2(n16344), .B1(n25254), .B2(n16342), .ZN(
        n24813) );
  NAND2_X2 U10468 ( .A1(n16344), .A2(n11634), .ZN(n16342) );
  NOR2_X2 U10470 ( .A1(n16346), .A2(n16347), .ZN(n16344) );
  NAND3_X2 U10472 ( .A1(n24833), .A2(n24832), .A3(n16218), .ZN(n12971) );
  NOR2_X2 U10473 ( .A1(n25249), .A2(n22385), .ZN(n16218) );
  OAI22_X2 U10480 ( .A1(n22385), .A2(n16353), .B1(n16348), .B2(n16354), .ZN(
        n24816) );
  OAI22_X2 U10483 ( .A1(n22386), .A2(n26292), .B1(n24833), .B2(n16348), .ZN(
        n24817) );
  NAND2_X2 U10484 ( .A1(n16347), .A2(n26292), .ZN(n16348) );
  NOR2_X2 U10485 ( .A1(n26293), .A2(n12844), .ZN(n16347) );
  NOR3_X2 U10486 ( .A1(n25400), .A2(n22386), .A3(n16298), .ZN(n12844) );
  NAND2_X2 U10487 ( .A1(n22384), .A2(n25249), .ZN(n16298) );
  OAI22_X2 U10494 ( .A1(n28822), .A2(n26293), .B1(n26305), .B2(n16358), .ZN(
        n24819) );
  OAI22_X2 U10497 ( .A1(n11788), .A2(n16358), .B1(n22422), .B2(n16360), .ZN(
        n24820) );
  NAND2_X2 U10506 ( .A1(n16364), .A2(n11634), .ZN(n16358) );
  NOR2_X2 U10509 ( .A1(n26135), .A2(n26293), .ZN(n16346) );
  NOR3_X2 U10513 ( .A1(n22423), .A2(n22422), .A3(n22424), .ZN(n16359) );
  NAND2_X2 U10519 ( .A1(n11876), .A2(n24894), .ZN(n13043) );
  NOR3_X2 U10521 ( .A1(n11878), .A2(n22420), .A3(n26129), .ZN(n11876) );
  NAND2_X2 U10523 ( .A1(n11220), .A2(n11200), .ZN(n11878) );
  NOR2_X2 U10526 ( .A1(n22419), .A2(n22418), .ZN(n11203) );
  NOR2_X2 U10527 ( .A1(n22415), .A2(n22414), .ZN(n11257) );
  DFF_X2 mac_b_reg_3_ ( .D(n25768), .CK(clk), .Q(n25769), .QN(n18903) );
  DFF_X2 mac_a3_reg_3_ ( .D(n23503), .CK(clk), .Q(n25739), .QN(n16855) );
  DFF_X2 mac_b_reg_2_ ( .D(n23101), .CK(clk), .Q(n4890), .QN(n18866) );
  DFF_X2 mac_b_reg_6_ ( .D(n23097), .CK(clk), .QN(n19014) );
  DFF_X2 mac_a3_reg_7_ ( .D(n23507), .CK(clk), .QN(n16707) );
  DFF_X2 mac_z_reg_1_ ( .D(n20554), .CK(clk), .Q(n25757), .QN(n20457) );
  DFF_X2 mac_a3_reg_4_ ( .D(n23504), .CK(clk), .QN(n16818) );
  DFF_X2 m_reg_5_ ( .D(n20561), .CK(clk), .QN(n20529) );
  DFF_X2 m_reg_2_ ( .D(n20558), .CK(clk), .QN(n20526) );
  DFF_X2 m_reg_1_ ( .D(n20557), .CK(clk), .Q(n25755), .QN(n20525) );
  DFF_X2 m_reg_6_ ( .D(n20562), .CK(clk), .Q(n5047), .QN(n20530) );
  DFF_X2 mac_b_reg_1_ ( .D(n25771), .CK(clk), .Q(n25772), .QN(n25984) );
  DFF_X2 m_reg_3_ ( .D(n20559), .CK(clk), .Q(n25779), .QN(n25778) );
  DFF_X2 mac_z_reg_7_ ( .D(n20548), .CK(clk), .Q(n643), .QN(n20067) );
  DFF_X2 mac_z_reg_2_ ( .D(n20553), .CK(clk), .QN(n20392) );
  DFF_X2 mac_z_reg_4_ ( .D(n20551), .CK(clk), .QN(n20262) );
  DFF_X2 dut__xxx__finish_reg ( .D(n22382), .CK(clk), .Q(dut__xxx__finish), 
        .QN(n16365) );
  DFF_X2 dut__dim__address_reg_7_ ( .D(n24649), .CK(clk), .Q(
        dut__dim__address[7]), .QN(n16366) );
  DFF_X2 dut__bvm__address_reg_1_ ( .D(n23265), .CK(clk), .Q(
        dut__bvm__address[1]), .QN(n18754) );
  DFF_X2 dut__dim__address_reg_2_ ( .D(n21420), .CK(clk), .Q(
        dut__dim__address[2]), .QN(n16371) );
  DFF_X2 dut__bvm__address_reg_3_ ( .D(n23267), .CK(clk), .Q(
        dut__bvm__address[3]), .QN(n18752) );
  DFF_X2 dut__bvm__address_reg_4_ ( .D(n23268), .CK(clk), .Q(
        dut__bvm__address[4]), .QN(n18751) );
  DFF_X2 dut__bvm__address_reg_5_ ( .D(n23269), .CK(clk), .Q(
        dut__bvm__address[5]), .QN(n18750) );
  DFF_X2 dut__dim__address_reg_0_ ( .D(n24644), .CK(clk), .Q(
        dut__dim__address[0]), .QN(n16373) );
  DFF_X2 dut__dim__address_reg_5_ ( .D(n24648), .CK(clk), .Q(
        dut__dim__address[5]), .QN(n16368) );
  DFF_X2 dut__bvm__address_reg_0_ ( .D(n23264), .CK(clk), .Q(
        dut__bvm__address[0]), .QN(n18755) );
  DFF_X2 dut__bvm__address_reg_2_ ( .D(n23266), .CK(clk), .Q(
        dut__bvm__address[2]), .QN(n18753) );
  DFF_X2 dut__dom__address_reg_0_ ( .D(n22428), .CK(clk), .Q(
        dut__dom__address[0]), .QN(n19482) );
  DFF_X2 dut__dom__address_reg_1_ ( .D(n22429), .CK(clk), .Q(
        dut__dom__address[1]), .QN(n19481) );
  DFF_X2 dut__dom__address_reg_2_ ( .D(n22430), .CK(clk), .Q(
        dut__dom__address[2]), .QN(n19480) );
  DFF_X2 dut__dom__enable_reg ( .D(n21151), .CK(clk), .Q(dut__dom__enable), 
        .QN(n19351) );
  DFF_X2 dut__dom__write_reg ( .D(n21150), .CK(clk), .Q(dut__dom__write), .QN(
        n19350) );
  DFF_X2 dut__bvm__address_reg_7_ ( .D(n21152), .CK(clk), .Q(
        dut__bvm__address[7]), .QN(n18748) );
  DFF_X2 dut__bvm__address_reg_8_ ( .D(n21153), .CK(clk), .Q(
        dut__bvm__address[8]), .QN(n18747) );
  DFF_X2 dut__bvm__address_reg_9_ ( .D(n21154), .CK(clk), .Q(
        dut__bvm__address[9]), .QN(n18746) );
  DFF_X2 dut__dim__address_reg_6_ ( .D(n21419), .CK(clk), .Q(
        dut__dim__address[6]), .QN(n16367) );
  DFF_X2 dut__dim__address_reg_4_ ( .D(n24647), .CK(clk), .Q(
        dut__dim__address[4]), .QN(n16369) );
  DFF_X2 dut__dim__address_reg_1_ ( .D(n24645), .CK(clk), .Q(
        dut__dim__address[1]), .QN(n16372) );
  DFF_X2 mac_a3_reg_5_ ( .D(n23505), .CK(clk), .Q(n25735), .QN(n16781) );
  DFF_X2 dut__dim__address_reg_3_ ( .D(n24646), .CK(clk), .Q(
        dut__dim__address[3]), .QN(n16370) );
  DFF_X2 mac_z_reg_5_ ( .D(n20550), .CK(clk), .Q(n25743), .QN(n20197) );
  DFF_X2 mac_z_reg_3_ ( .D(n20552), .CK(clk), .Q(n25749), .QN(n20327) );
  DFF_X2 mac_a3_reg_1_ ( .D(n23501), .CK(clk), .Q(n25745), .QN(n16929) );
  DFF_X2 mac_b_reg_0_ ( .D(n23103), .CK(clk), .Q(n4888), .QN(n18792) );
  DFF_X2 m_reg_7_ ( .D(n20563), .CK(clk), .Q(n5048), .QN(n20531) );
  DFF_X2 mac_a3_reg_0_ ( .D(n23500), .CK(clk), .QN(n16966) );
  DFF_X2 m_reg_4_ ( .D(n20560), .CK(clk), .QN(n20528) );
  DFF_X2 mac_b_reg_4_ ( .D(n23099), .CK(clk), .QN(n18940) );
  DFF_X2 mac_a3_reg_2_ ( .D(n23502), .CK(clk), .Q(n4906), .QN(n16892) );
  DFF_X2 dut__bvm__enable_reg ( .D(n22447), .CK(clk), .Q(dut__bvm__enable) );
  DFF_X2 z_reg_62__15_ ( .D(n25399), .CK(clk), .Q(n26153), .QN(n28694) );
  DFF_X2 z_reg_57__15_ ( .D(n25398), .CK(clk), .Q(n26167), .QN(n28510) );
  DFF_X2 z_reg_52__15_ ( .D(n25397), .CK(clk), .Q(n26141), .QN(n28256) );
  DFF_X2 z_reg_49__15_ ( .D(n25396), .CK(clk), .Q(n26140), .QN(n28257) );
  DFF_X2 z_reg_14__15_ ( .D(n25097), .CK(clk), .Q(n19513) );
  DFF_X2 z_reg_11__15_ ( .D(n25395), .CK(clk), .Q(n26152), .QN(n28695) );
  DFF_X2 z_reg_6__15_ ( .D(n25394), .CK(clk), .Q(n26181), .QN(n28381) );
  DFF_X2 z_reg_3__15_ ( .D(n25103), .CK(clk), .Q(n19508) );
  DFF_X2 z_reg_28__15_ ( .D(n25393), .CK(clk), .Q(n26168), .QN(n28509) );
  DFF_X2 z_reg_25__15_ ( .D(n25091), .CK(clk), .Q(n19504) );
  DFF_X2 z_reg_20__15_ ( .D(n25392), .CK(clk), .Q(n26142), .QN(n28255) );
  DFF_X2 z_reg_17__15_ ( .D(n25090), .CK(clk), .Q(n19500) );
  DFF_X2 z_reg_46__15_ ( .D(n25391), .CK(clk), .Q(n26154), .QN(n28693) );
  DFF_X2 z_reg_43__15_ ( .D(n25095), .CK(clk), .Q(n19496) );
  DFF_X2 z_reg_38__15_ ( .D(n25390), .CK(clk), .Q(n26182), .QN(n28380) );
  DFF_X2 z_reg_35__15_ ( .D(n25094), .CK(clk), .Q(n19492) );
  DFF_X2 z_reg_48__15_ ( .D(n25101), .CK(clk), .Q(n19483) );
  DFF_X2 z_reg_63__15_ ( .D(n25093), .CK(clk), .Q(n19490) );
  DFF_X2 z_reg_53__15_ ( .D(n25092), .CK(clk), .Q(n19486) );
  DFF_X2 z_reg_24__15_ ( .D(n25089), .CK(clk), .Q(n19503) );
  DFF_X2 z_reg_16__15_ ( .D(n25088), .CK(clk), .Q(n19499) );
  DFF_X2 z_reg_42__15_ ( .D(n25087), .CK(clk), .Q(n19495) );
  DFF_X2 z_reg_34__15_ ( .D(n25086), .CK(clk), .Q(n19491) );
  DFF_X2 z_reg_47__15_ ( .D(n25389), .CK(clk), .Q(n26155), .QN(n28692) );
  DFF_X2 z_reg_39__15_ ( .D(n25388), .CK(clk), .Q(n26183), .QN(n28379) );
  DFF_X2 z_reg_29__15_ ( .D(n25387), .CK(clk), .Q(n26169), .QN(n28508) );
  DFF_X2 z_reg_21__15_ ( .D(n25386), .CK(clk), .Q(n26143), .QN(n28254) );
  DFF_X2 z_reg_15__15_ ( .D(n25102), .CK(clk), .Q(n19514) );
  DFF_X2 z_reg_7__15_ ( .D(n25385), .CK(clk), .Q(n26180), .QN(n28382) );
  DFF_X2 z_reg_10__15_ ( .D(n25361), .CK(clk), .Q(n26151), .QN(n28696) );
  DFF_X2 z_reg_2__15_ ( .D(n25083), .CK(clk), .Q(n19507) );
  DFF_X2 z_reg_56__15_ ( .D(n25081), .CK(clk), .Q(n19487) );
  DFF_X2 output_store_reg_5__15_ ( .D(n25261), .CK(clk), .Q(n26165), .QN(
        n28818) );
  DFF_X2 z_reg_62__14_ ( .D(n22942), .CK(clk), .QN(n28685) );
  DFF_X2 z_reg_62__13_ ( .D(n22952), .CK(clk), .QN(n28674) );
  DFF_X2 z_reg_62__12_ ( .D(n22962), .CK(clk), .QN(n28663) );
  DFF_X2 z_reg_62__11_ ( .D(n22972), .CK(clk), .QN(n28652) );
  DFF_X2 z_reg_62__10_ ( .D(n22982), .CK(clk), .QN(n28641) );
  DFF_X2 z_reg_62__9_ ( .D(n22992), .CK(clk), .QN(n28630) );
  DFF_X2 z_reg_62__8_ ( .D(n23002), .CK(clk), .QN(n28619) );
  DFF_X2 z_reg_62__7_ ( .D(n23012), .CK(clk), .QN(n28608) );
  DFF_X2 z_reg_62__6_ ( .D(n23022), .CK(clk), .QN(n28597) );
  DFF_X2 z_reg_62__5_ ( .D(n23032), .CK(clk), .QN(n28586) );
  DFF_X2 z_reg_62__4_ ( .D(n23042), .CK(clk), .QN(n28575) );
  DFF_X2 z_reg_62__3_ ( .D(n23052), .CK(clk), .QN(n28560) );
  DFF_X2 z_reg_62__2_ ( .D(n23062), .CK(clk), .QN(n28545) );
  DFF_X2 z_reg_62__1_ ( .D(n23072), .CK(clk), .QN(n28530) );
  DFF_X2 z_reg_62__0_ ( .D(n23082), .CK(clk), .QN(n28515) );
  DFF_X2 z_reg_57__14_ ( .D(n22842), .CK(clk), .QN(n28505) );
  DFF_X2 z_reg_57__13_ ( .D(n22848), .CK(clk), .QN(n28498) );
  DFF_X2 z_reg_57__12_ ( .D(n22854), .CK(clk), .QN(n28491) );
  DFF_X2 z_reg_57__11_ ( .D(n22860), .CK(clk), .QN(n28484) );
  DFF_X2 z_reg_57__10_ ( .D(n22866), .CK(clk), .QN(n28477) );
  DFF_X2 z_reg_57__9_ ( .D(n22872), .CK(clk), .QN(n28470) );
  DFF_X2 z_reg_57__8_ ( .D(n22878), .CK(clk), .QN(n28463) );
  DFF_X2 z_reg_57__7_ ( .D(n22884), .CK(clk), .QN(n28456) );
  DFF_X2 z_reg_57__6_ ( .D(n22890), .CK(clk), .QN(n28449) );
  DFF_X2 z_reg_57__5_ ( .D(n22896), .CK(clk), .QN(n28442) );
  DFF_X2 z_reg_57__4_ ( .D(n22902), .CK(clk), .QN(n28435) );
  DFF_X2 z_reg_57__3_ ( .D(n22908), .CK(clk), .QN(n28423) );
  DFF_X2 z_reg_57__2_ ( .D(n22914), .CK(clk), .QN(n28411) );
  DFF_X2 z_reg_57__1_ ( .D(n22920), .CK(clk), .QN(n28399) );
  DFF_X2 z_reg_57__0_ ( .D(n22926), .CK(clk), .QN(n28387) );
  DFF_X2 z_reg_52__8_ ( .D(n22636), .CK(clk), .QN(n28202) );
  DFF_X2 z_reg_52__7_ ( .D(n22644), .CK(clk), .QN(n28194) );
  DFF_X2 z_reg_52__6_ ( .D(n22652), .CK(clk), .QN(n28186) );
  DFF_X2 z_reg_52__5_ ( .D(n22660), .CK(clk), .QN(n28178) );
  DFF_X2 z_reg_52__4_ ( .D(n22668), .CK(clk), .QN(n28170) );
  DFF_X2 z_reg_52__3_ ( .D(n22676), .CK(clk), .QN(n28162) );
  DFF_X2 z_reg_52__2_ ( .D(n22684), .CK(clk), .QN(n28154) );
  DFF_X2 z_reg_52__1_ ( .D(n22692), .CK(clk), .QN(n28146) );
  DFF_X2 z_reg_52__0_ ( .D(n22700), .CK(clk), .QN(n28138) );
  DFF_X2 z_reg_49__8_ ( .D(n22637), .CK(clk), .QN(n28203) );
  DFF_X2 z_reg_49__7_ ( .D(n22645), .CK(clk), .QN(n28195) );
  DFF_X2 z_reg_49__6_ ( .D(n22653), .CK(clk), .QN(n28187) );
  DFF_X2 z_reg_49__5_ ( .D(n22661), .CK(clk), .QN(n28179) );
  DFF_X2 z_reg_49__4_ ( .D(n22669), .CK(clk), .QN(n28171) );
  DFF_X2 z_reg_49__3_ ( .D(n22677), .CK(clk), .QN(n28163) );
  DFF_X2 z_reg_49__2_ ( .D(n22685), .CK(clk), .QN(n28155) );
  DFF_X2 z_reg_49__1_ ( .D(n22693), .CK(clk), .QN(n28147) );
  DFF_X2 z_reg_49__0_ ( .D(n22701), .CK(clk), .QN(n28139) );
  DFF_X2 z_reg_14__14_ ( .D(n22943), .CK(clk), .Q(n19578), .QN(n28686) );
  DFF_X2 z_reg_14__13_ ( .D(n22953), .CK(clk), .Q(n19643), .QN(n28675) );
  DFF_X2 z_reg_14__12_ ( .D(n22963), .CK(clk), .Q(n19708), .QN(n28664) );
  DFF_X2 z_reg_14__11_ ( .D(n22973), .CK(clk), .Q(n19773), .QN(n28653) );
  DFF_X2 z_reg_14__10_ ( .D(n22983), .CK(clk), .Q(n19838), .QN(n28642) );
  DFF_X2 z_reg_14__9_ ( .D(n22993), .CK(clk), .Q(n19903), .QN(n28631) );
  DFF_X2 z_reg_14__8_ ( .D(n23003), .CK(clk), .Q(n19968), .QN(n28620) );
  DFF_X2 z_reg_14__7_ ( .D(n23013), .CK(clk), .Q(n20033), .QN(n28609) );
  DFF_X2 z_reg_14__6_ ( .D(n23023), .CK(clk), .Q(n20098), .QN(n28598) );
  DFF_X2 z_reg_14__5_ ( .D(n23033), .CK(clk), .Q(n20163), .QN(n28587) );
  DFF_X2 z_reg_14__4_ ( .D(n23043), .CK(clk), .Q(n20228), .QN(n28576) );
  DFF_X2 z_reg_14__3_ ( .D(n23053), .CK(clk), .Q(n20293), .QN(n28561) );
  DFF_X2 z_reg_14__2_ ( .D(n23063), .CK(clk), .Q(n20358), .QN(n28546) );
  DFF_X2 z_reg_14__1_ ( .D(n23073), .CK(clk), .Q(n20423), .QN(n28531) );
  DFF_X2 z_reg_14__0_ ( .D(n23083), .CK(clk), .Q(n20489), .QN(n28516) );
  DFF_X2 z_reg_11__14_ ( .D(n22944), .CK(clk), .QN(n28687) );
  DFF_X2 z_reg_11__13_ ( .D(n22954), .CK(clk), .QN(n28676) );
  DFF_X2 z_reg_11__12_ ( .D(n22964), .CK(clk), .QN(n28665) );
  DFF_X2 z_reg_11__11_ ( .D(n22974), .CK(clk), .QN(n28654) );
  DFF_X2 z_reg_11__10_ ( .D(n22984), .CK(clk), .QN(n28643) );
  DFF_X2 z_reg_11__9_ ( .D(n22994), .CK(clk), .QN(n28632) );
  DFF_X2 z_reg_11__8_ ( .D(n23004), .CK(clk), .QN(n28621) );
  DFF_X2 z_reg_11__7_ ( .D(n23014), .CK(clk), .QN(n28610) );
  DFF_X2 z_reg_11__6_ ( .D(n23024), .CK(clk), .QN(n28599) );
  DFF_X2 z_reg_11__5_ ( .D(n23034), .CK(clk), .QN(n28588) );
  DFF_X2 z_reg_11__4_ ( .D(n23044), .CK(clk), .QN(n28577) );
  DFF_X2 z_reg_11__3_ ( .D(n23054), .CK(clk), .QN(n28562) );
  DFF_X2 z_reg_11__2_ ( .D(n23064), .CK(clk), .QN(n28547) );
  DFF_X2 z_reg_11__1_ ( .D(n23074), .CK(clk), .QN(n28532) );
  DFF_X2 z_reg_11__0_ ( .D(n23084), .CK(clk), .QN(n28517) );
  DFF_X2 z_reg_6__8_ ( .D(n22764), .CK(clk), .QN(n28326) );
  DFF_X2 z_reg_6__7_ ( .D(n22772), .CK(clk), .QN(n28318) );
  DFF_X2 z_reg_6__6_ ( .D(n22780), .CK(clk), .QN(n28310) );
  DFF_X2 z_reg_6__5_ ( .D(n22788), .CK(clk), .QN(n28302) );
  DFF_X2 z_reg_6__4_ ( .D(n22796), .CK(clk), .QN(n28294) );
  DFF_X2 z_reg_6__3_ ( .D(n22804), .CK(clk), .QN(n28286) );
  DFF_X2 z_reg_6__2_ ( .D(n22812), .CK(clk), .QN(n28278) );
  DFF_X2 z_reg_6__1_ ( .D(n22820), .CK(clk), .QN(n28270) );
  DFF_X2 z_reg_6__0_ ( .D(n22828), .CK(clk), .QN(n28262) );
  DFF_X2 z_reg_3__8_ ( .D(n22765), .CK(clk), .Q(n19963), .QN(n28327) );
  DFF_X2 z_reg_3__7_ ( .D(n22773), .CK(clk), .Q(n20028), .QN(n28319) );
  DFF_X2 z_reg_3__6_ ( .D(n22781), .CK(clk), .Q(n20093), .QN(n28311) );
  DFF_X2 z_reg_3__5_ ( .D(n22789), .CK(clk), .Q(n20158), .QN(n28303) );
  DFF_X2 z_reg_3__4_ ( .D(n22797), .CK(clk), .Q(n20223), .QN(n28295) );
  DFF_X2 z_reg_3__3_ ( .D(n22805), .CK(clk), .Q(n20288), .QN(n28287) );
  DFF_X2 z_reg_3__2_ ( .D(n22813), .CK(clk), .Q(n20353), .QN(n28279) );
  DFF_X2 z_reg_3__1_ ( .D(n22821), .CK(clk), .Q(n20418), .QN(n28271) );
  DFF_X2 z_reg_3__0_ ( .D(n22829), .CK(clk), .Q(n20484), .QN(n28263) );
  DFF_X2 z_reg_46__14_ ( .D(n22939), .CK(clk), .QN(n28682) );
  DFF_X2 z_reg_46__13_ ( .D(n22949), .CK(clk), .QN(n28671) );
  DFF_X2 z_reg_46__12_ ( .D(n22959), .CK(clk), .QN(n28660) );
  DFF_X2 z_reg_46__11_ ( .D(n22969), .CK(clk), .QN(n28649) );
  DFF_X2 z_reg_46__10_ ( .D(n22979), .CK(clk), .QN(n28638) );
  DFF_X2 z_reg_46__9_ ( .D(n22989), .CK(clk), .QN(n28627) );
  DFF_X2 z_reg_46__8_ ( .D(n22999), .CK(clk), .QN(n28616) );
  DFF_X2 z_reg_46__7_ ( .D(n23009), .CK(clk), .QN(n28605) );
  DFF_X2 z_reg_46__6_ ( .D(n23019), .CK(clk), .QN(n28594) );
  DFF_X2 z_reg_46__5_ ( .D(n23029), .CK(clk), .QN(n28583) );
  DFF_X2 z_reg_46__4_ ( .D(n23039), .CK(clk), .QN(n28572) );
  DFF_X2 z_reg_46__3_ ( .D(n23049), .CK(clk), .QN(n28557) );
  DFF_X2 z_reg_46__2_ ( .D(n23059), .CK(clk), .QN(n28542) );
  DFF_X2 z_reg_46__1_ ( .D(n23069), .CK(clk), .QN(n28527) );
  DFF_X2 z_reg_46__0_ ( .D(n23079), .CK(clk), .QN(n28512) );
  DFF_X2 z_reg_43__14_ ( .D(n22940), .CK(clk), .Q(n19561), .QN(n28683) );
  DFF_X2 z_reg_43__13_ ( .D(n22950), .CK(clk), .Q(n19626), .QN(n28672) );
  DFF_X2 z_reg_43__12_ ( .D(n22960), .CK(clk), .Q(n19691), .QN(n28661) );
  DFF_X2 z_reg_43__11_ ( .D(n22970), .CK(clk), .Q(n19756), .QN(n28650) );
  DFF_X2 z_reg_43__10_ ( .D(n22980), .CK(clk), .Q(n19821), .QN(n28639) );
  DFF_X2 z_reg_43__9_ ( .D(n22990), .CK(clk), .Q(n19886), .QN(n28628) );
  DFF_X2 z_reg_43__8_ ( .D(n23000), .CK(clk), .Q(n19951), .QN(n28617) );
  DFF_X2 z_reg_43__7_ ( .D(n23010), .CK(clk), .Q(n20016), .QN(n28606) );
  DFF_X2 z_reg_43__6_ ( .D(n23020), .CK(clk), .Q(n20081), .QN(n28595) );
  DFF_X2 z_reg_43__5_ ( .D(n23030), .CK(clk), .Q(n20146), .QN(n28584) );
  DFF_X2 z_reg_43__4_ ( .D(n23040), .CK(clk), .Q(n20211), .QN(n28573) );
  DFF_X2 z_reg_43__3_ ( .D(n23050), .CK(clk), .Q(n20276), .QN(n28558) );
  DFF_X2 z_reg_43__2_ ( .D(n23060), .CK(clk), .Q(n20341), .QN(n28543) );
  DFF_X2 z_reg_43__1_ ( .D(n23070), .CK(clk), .Q(n20406), .QN(n28528) );
  DFF_X2 z_reg_43__0_ ( .D(n23080), .CK(clk), .Q(n20472), .QN(n28513) );
  DFF_X2 z_reg_38__8_ ( .D(n22761), .CK(clk), .QN(n28323) );
  DFF_X2 z_reg_38__7_ ( .D(n22769), .CK(clk), .QN(n28315) );
  DFF_X2 z_reg_38__6_ ( .D(n22777), .CK(clk), .QN(n28307) );
  DFF_X2 z_reg_38__5_ ( .D(n22785), .CK(clk), .QN(n28299) );
  DFF_X2 z_reg_38__4_ ( .D(n22793), .CK(clk), .QN(n28291) );
  DFF_X2 z_reg_38__3_ ( .D(n22801), .CK(clk), .QN(n28283) );
  DFF_X2 z_reg_38__2_ ( .D(n22809), .CK(clk), .QN(n28275) );
  DFF_X2 z_reg_38__1_ ( .D(n22817), .CK(clk), .QN(n28267) );
  DFF_X2 z_reg_38__0_ ( .D(n22825), .CK(clk), .QN(n28259) );
  DFF_X2 z_reg_35__8_ ( .D(n22762), .CK(clk), .Q(n19947), .QN(n28324) );
  DFF_X2 z_reg_35__7_ ( .D(n22770), .CK(clk), .Q(n20012), .QN(n28316) );
  DFF_X2 z_reg_35__6_ ( .D(n22778), .CK(clk), .Q(n20077), .QN(n28308) );
  DFF_X2 z_reg_35__5_ ( .D(n22786), .CK(clk), .Q(n20142), .QN(n28300) );
  DFF_X2 z_reg_35__4_ ( .D(n22794), .CK(clk), .Q(n20207), .QN(n28292) );
  DFF_X2 z_reg_35__3_ ( .D(n22802), .CK(clk), .Q(n20272), .QN(n28284) );
  DFF_X2 z_reg_35__2_ ( .D(n22810), .CK(clk), .Q(n20337), .QN(n28276) );
  DFF_X2 z_reg_35__1_ ( .D(n22818), .CK(clk), .Q(n20402), .QN(n28268) );
  DFF_X2 z_reg_35__0_ ( .D(n22826), .CK(clk), .Q(n20468), .QN(n28260) );
  DFF_X2 z_reg_28__14_ ( .D(n22839), .CK(clk), .QN(n28502) );
  DFF_X2 z_reg_28__13_ ( .D(n22845), .CK(clk), .QN(n28495) );
  DFF_X2 z_reg_28__12_ ( .D(n22851), .CK(clk), .QN(n28488) );
  DFF_X2 z_reg_28__11_ ( .D(n22857), .CK(clk), .QN(n28481) );
  DFF_X2 z_reg_28__10_ ( .D(n22863), .CK(clk), .QN(n28474) );
  DFF_X2 z_reg_28__9_ ( .D(n22869), .CK(clk), .QN(n28467) );
  DFF_X2 z_reg_28__8_ ( .D(n22875), .CK(clk), .QN(n28460) );
  DFF_X2 z_reg_28__7_ ( .D(n22881), .CK(clk), .QN(n28453) );
  DFF_X2 z_reg_28__6_ ( .D(n22887), .CK(clk), .QN(n28446) );
  DFF_X2 z_reg_28__5_ ( .D(n22893), .CK(clk), .QN(n28439) );
  DFF_X2 z_reg_28__4_ ( .D(n22899), .CK(clk), .QN(n28432) );
  DFF_X2 z_reg_28__3_ ( .D(n22905), .CK(clk), .QN(n28420) );
  DFF_X2 z_reg_28__2_ ( .D(n22911), .CK(clk), .QN(n28408) );
  DFF_X2 z_reg_28__1_ ( .D(n22917), .CK(clk), .QN(n28396) );
  DFF_X2 z_reg_28__0_ ( .D(n22923), .CK(clk), .QN(n28384) );
  DFF_X2 z_reg_25__14_ ( .D(n22840), .CK(clk), .Q(n19569), .QN(n28503) );
  DFF_X2 z_reg_25__13_ ( .D(n22846), .CK(clk), .Q(n19634), .QN(n28496) );
  DFF_X2 z_reg_25__12_ ( .D(n22852), .CK(clk), .Q(n19699), .QN(n28489) );
  DFF_X2 z_reg_25__11_ ( .D(n22858), .CK(clk), .Q(n19764), .QN(n28482) );
  DFF_X2 z_reg_25__10_ ( .D(n22864), .CK(clk), .Q(n19829), .QN(n28475) );
  DFF_X2 z_reg_25__9_ ( .D(n22870), .CK(clk), .Q(n19894), .QN(n28468) );
  DFF_X2 z_reg_25__8_ ( .D(n22876), .CK(clk), .Q(n19959), .QN(n28461) );
  DFF_X2 z_reg_25__7_ ( .D(n22882), .CK(clk), .Q(n20024), .QN(n28454) );
  DFF_X2 z_reg_25__6_ ( .D(n22888), .CK(clk), .Q(n20089), .QN(n28447) );
  DFF_X2 z_reg_25__5_ ( .D(n22894), .CK(clk), .Q(n20154), .QN(n28440) );
  DFF_X2 z_reg_25__4_ ( .D(n22900), .CK(clk), .Q(n20219), .QN(n28433) );
  DFF_X2 z_reg_25__3_ ( .D(n22906), .CK(clk), .Q(n20284), .QN(n28421) );
  DFF_X2 z_reg_25__2_ ( .D(n22912), .CK(clk), .Q(n20349), .QN(n28409) );
  DFF_X2 z_reg_25__1_ ( .D(n22918), .CK(clk), .Q(n20414), .QN(n28397) );
  DFF_X2 z_reg_25__0_ ( .D(n22924), .CK(clk), .Q(n20480), .QN(n28385) );
  DFF_X2 z_reg_20__8_ ( .D(n22633), .CK(clk), .QN(n28199) );
  DFF_X2 z_reg_20__7_ ( .D(n22641), .CK(clk), .QN(n28191) );
  DFF_X2 z_reg_20__6_ ( .D(n22649), .CK(clk), .QN(n28183) );
  DFF_X2 z_reg_20__5_ ( .D(n22657), .CK(clk), .QN(n28175) );
  DFF_X2 z_reg_20__4_ ( .D(n22665), .CK(clk), .QN(n28167) );
  DFF_X2 z_reg_20__3_ ( .D(n22673), .CK(clk), .QN(n28159) );
  DFF_X2 z_reg_20__2_ ( .D(n22681), .CK(clk), .QN(n28151) );
  DFF_X2 z_reg_20__1_ ( .D(n22689), .CK(clk), .QN(n28143) );
  DFF_X2 z_reg_20__0_ ( .D(n22697), .CK(clk), .QN(n28135) );
  DFF_X2 z_reg_17__8_ ( .D(n22634), .CK(clk), .Q(n19955), .QN(n28200) );
  DFF_X2 z_reg_17__7_ ( .D(n22642), .CK(clk), .Q(n20020), .QN(n28192) );
  DFF_X2 z_reg_17__6_ ( .D(n22650), .CK(clk), .Q(n20085), .QN(n28184) );
  DFF_X2 z_reg_17__5_ ( .D(n22658), .CK(clk), .Q(n20150), .QN(n28176) );
  DFF_X2 z_reg_17__4_ ( .D(n22666), .CK(clk), .Q(n20215), .QN(n28168) );
  DFF_X2 z_reg_17__3_ ( .D(n22674), .CK(clk), .Q(n20280), .QN(n28160) );
  DFF_X2 z_reg_17__2_ ( .D(n22682), .CK(clk), .Q(n20345), .QN(n28152) );
  DFF_X2 z_reg_17__1_ ( .D(n22690), .CK(clk), .Q(n20410), .QN(n28144) );
  DFF_X2 z_reg_17__0_ ( .D(n22698), .CK(clk), .Q(n20476), .QN(n28136) );
  DFF_X2 flag_zsynch_reg ( .D(n23440), .CK(clk), .Q(n20458), .QN(n27805) );
  DFF_X2 z_reg_10__14_ ( .D(n22946), .CK(clk), .QN(n28689) );
  DFF_X2 z_reg_10__13_ ( .D(n22956), .CK(clk), .QN(n28678) );
  DFF_X2 z_reg_10__11_ ( .D(n22976), .CK(clk), .QN(n28656) );
  DFF_X2 z_reg_10__10_ ( .D(n22986), .CK(clk), .QN(n28645) );
  DFF_X2 z_reg_10__8_ ( .D(n23006), .CK(clk), .QN(n28623) );
  DFF_X2 z_reg_10__4_ ( .D(n23046), .CK(clk), .QN(n28579) );
  DFF_X2 z_reg_10__2_ ( .D(n23066), .CK(clk), .QN(n28549) );
  DFF_X2 z_reg_10__0_ ( .D(n23086), .CK(clk), .QN(n28519) );
  DFF_X2 z_reg_56__14_ ( .D(n22843), .CK(clk), .Q(n19552), .QN(n28506) );
  DFF_X2 z_reg_56__13_ ( .D(n22849), .CK(clk), .Q(n19617), .QN(n28499) );
  DFF_X2 z_reg_56__12_ ( .D(n22855), .CK(clk), .Q(n19682), .QN(n28492) );
  DFF_X2 z_reg_56__11_ ( .D(n22861), .CK(clk), .Q(n19747), .QN(n28485) );
  DFF_X2 z_reg_56__10_ ( .D(n22867), .CK(clk), .Q(n19812), .QN(n28478) );
  DFF_X2 z_reg_56__9_ ( .D(n22873), .CK(clk), .Q(n19877), .QN(n28471) );
  DFF_X2 z_reg_56__8_ ( .D(n22879), .CK(clk), .Q(n19942), .QN(n28464) );
  DFF_X2 z_reg_56__7_ ( .D(n22885), .CK(clk), .Q(n20007), .QN(n28457) );
  DFF_X2 z_reg_56__6_ ( .D(n22891), .CK(clk), .Q(n20072), .QN(n28450) );
  DFF_X2 z_reg_56__5_ ( .D(n22897), .CK(clk), .Q(n20137), .QN(n28443) );
  DFF_X2 z_reg_56__4_ ( .D(n22903), .CK(clk), .Q(n20202), .QN(n28436) );
  DFF_X2 z_reg_56__3_ ( .D(n22909), .CK(clk), .Q(n20267), .QN(n28424) );
  DFF_X2 z_reg_56__2_ ( .D(n22915), .CK(clk), .Q(n20332), .QN(n28412) );
  DFF_X2 z_reg_56__1_ ( .D(n22921), .CK(clk), .Q(n20397), .QN(n28400) );
  DFF_X2 z_reg_56__0_ ( .D(n22927), .CK(clk), .Q(n20463), .QN(n28388) );
  DFF_X2 z_reg_48__8_ ( .D(n22638), .CK(clk), .Q(n19938), .QN(n28204) );
  DFF_X2 z_reg_48__7_ ( .D(n22646), .CK(clk), .Q(n20003), .QN(n28196) );
  DFF_X2 z_reg_48__6_ ( .D(n22654), .CK(clk), .Q(n20068), .QN(n28188) );
  DFF_X2 z_reg_48__5_ ( .D(n22662), .CK(clk), .Q(n20133), .QN(n28180) );
  DFF_X2 z_reg_48__4_ ( .D(n22670), .CK(clk), .Q(n20198), .QN(n28172) );
  DFF_X2 z_reg_48__3_ ( .D(n22678), .CK(clk), .Q(n20263), .QN(n28164) );
  DFF_X2 z_reg_48__2_ ( .D(n22686), .CK(clk), .Q(n20328), .QN(n28156) );
  DFF_X2 z_reg_48__1_ ( .D(n22694), .CK(clk), .Q(n20393), .QN(n28148) );
  DFF_X2 z_reg_48__0_ ( .D(n22702), .CK(clk), .Q(n20459), .QN(n28140) );
  DFF_X2 z_reg_2__8_ ( .D(n22767), .CK(clk), .Q(n19962), .QN(n28329) );
  DFF_X2 z_reg_2__5_ ( .D(n22791), .CK(clk), .Q(n20157), .QN(n28305) );
  DFF_X2 z_reg_2__3_ ( .D(n22807), .CK(clk), .Q(n20287), .QN(n28289) );
  DFF_X2 z_reg_2__2_ ( .D(n22815), .CK(clk), .Q(n20352), .QN(n28281) );
  DFF_X2 z_reg_2__1_ ( .D(n22823), .CK(clk), .Q(n20417), .QN(n28273) );
  DFF_X2 z_reg_2__0_ ( .D(n22831), .CK(clk), .Q(n20483), .QN(n28265) );
  DFF_X2 z_reg_10__12_ ( .D(n22966), .CK(clk), .QN(n28667) );
  DFF_X2 z_reg_10__9_ ( .D(n22996), .CK(clk), .QN(n28634) );
  DFF_X2 z_reg_10__7_ ( .D(n23016), .CK(clk), .QN(n28612) );
  DFF_X2 z_reg_10__6_ ( .D(n23026), .CK(clk), .QN(n28601) );
  DFF_X2 z_reg_10__5_ ( .D(n23036), .CK(clk), .QN(n28590) );
  DFF_X2 z_reg_10__3_ ( .D(n23056), .CK(clk), .QN(n28564) );
  DFF_X2 z_reg_10__1_ ( .D(n23076), .CK(clk), .QN(n28534) );
  DFF_X2 z_reg_52__14_ ( .D(n22588), .CK(clk), .QN(n28250) );
  DFF_X2 z_reg_52__13_ ( .D(n22596), .CK(clk), .QN(n28242) );
  DFF_X2 z_reg_52__12_ ( .D(n22604), .CK(clk), .QN(n28234) );
  DFF_X2 z_reg_52__11_ ( .D(n22612), .CK(clk), .QN(n28226) );
  DFF_X2 z_reg_52__10_ ( .D(n22620), .CK(clk), .QN(n28218) );
  DFF_X2 z_reg_52__9_ ( .D(n22628), .CK(clk), .QN(n28210) );
  DFF_X2 z_reg_49__14_ ( .D(n22589), .CK(clk), .QN(n28251) );
  DFF_X2 z_reg_49__13_ ( .D(n22597), .CK(clk), .QN(n28243) );
  DFF_X2 z_reg_49__12_ ( .D(n22605), .CK(clk), .QN(n28235) );
  DFF_X2 z_reg_49__11_ ( .D(n22613), .CK(clk), .QN(n28227) );
  DFF_X2 z_reg_49__10_ ( .D(n22621), .CK(clk), .QN(n28219) );
  DFF_X2 z_reg_49__9_ ( .D(n22629), .CK(clk), .QN(n28211) );
  DFF_X2 z_reg_6__14_ ( .D(n22716), .CK(clk), .QN(n28374) );
  DFF_X2 z_reg_6__13_ ( .D(n22724), .CK(clk), .QN(n28366) );
  DFF_X2 z_reg_6__12_ ( .D(n22732), .CK(clk), .QN(n28358) );
  DFF_X2 z_reg_6__11_ ( .D(n22740), .CK(clk), .QN(n28350) );
  DFF_X2 z_reg_6__10_ ( .D(n22748), .CK(clk), .QN(n28342) );
  DFF_X2 z_reg_6__9_ ( .D(n22756), .CK(clk), .QN(n28334) );
  DFF_X2 z_reg_3__14_ ( .D(n22717), .CK(clk), .Q(n19573), .QN(n28375) );
  DFF_X2 z_reg_3__13_ ( .D(n22725), .CK(clk), .Q(n19638), .QN(n28367) );
  DFF_X2 z_reg_3__12_ ( .D(n22733), .CK(clk), .Q(n19703), .QN(n28359) );
  DFF_X2 z_reg_3__11_ ( .D(n22741), .CK(clk), .Q(n19768), .QN(n28351) );
  DFF_X2 z_reg_3__10_ ( .D(n22749), .CK(clk), .Q(n19833), .QN(n28343) );
  DFF_X2 z_reg_3__9_ ( .D(n22757), .CK(clk), .Q(n19898), .QN(n28335) );
  DFF_X2 z_reg_20__14_ ( .D(n22585), .CK(clk), .QN(n28247) );
  DFF_X2 z_reg_20__13_ ( .D(n22593), .CK(clk), .QN(n28239) );
  DFF_X2 z_reg_20__12_ ( .D(n22601), .CK(clk), .QN(n28231) );
  DFF_X2 z_reg_20__11_ ( .D(n22609), .CK(clk), .QN(n28223) );
  DFF_X2 z_reg_20__10_ ( .D(n22617), .CK(clk), .QN(n28215) );
  DFF_X2 z_reg_20__9_ ( .D(n22625), .CK(clk), .QN(n28207) );
  DFF_X2 z_reg_17__14_ ( .D(n22586), .CK(clk), .Q(n19565), .QN(n28248) );
  DFF_X2 z_reg_17__13_ ( .D(n22594), .CK(clk), .Q(n19630), .QN(n28240) );
  DFF_X2 z_reg_17__12_ ( .D(n22602), .CK(clk), .Q(n19695), .QN(n28232) );
  DFF_X2 z_reg_17__11_ ( .D(n22610), .CK(clk), .Q(n19760), .QN(n28224) );
  DFF_X2 z_reg_17__10_ ( .D(n22618), .CK(clk), .Q(n19825), .QN(n28216) );
  DFF_X2 z_reg_17__9_ ( .D(n22626), .CK(clk), .Q(n19890), .QN(n28208) );
  DFF_X2 z_reg_38__14_ ( .D(n22713), .CK(clk), .QN(n28371) );
  DFF_X2 z_reg_38__13_ ( .D(n22721), .CK(clk), .QN(n28363) );
  DFF_X2 z_reg_38__12_ ( .D(n22729), .CK(clk), .QN(n28355) );
  DFF_X2 z_reg_38__11_ ( .D(n22737), .CK(clk), .QN(n28347) );
  DFF_X2 z_reg_38__10_ ( .D(n22745), .CK(clk), .QN(n28339) );
  DFF_X2 z_reg_38__9_ ( .D(n22753), .CK(clk), .QN(n28331) );
  DFF_X2 z_reg_35__14_ ( .D(n22714), .CK(clk), .Q(n19557), .QN(n28372) );
  DFF_X2 z_reg_35__13_ ( .D(n22722), .CK(clk), .Q(n19622), .QN(n28364) );
  DFF_X2 z_reg_35__12_ ( .D(n22730), .CK(clk), .Q(n19687), .QN(n28356) );
  DFF_X2 z_reg_35__11_ ( .D(n22738), .CK(clk), .Q(n19752), .QN(n28348) );
  DFF_X2 z_reg_35__10_ ( .D(n22746), .CK(clk), .Q(n19817), .QN(n28340) );
  DFF_X2 z_reg_35__9_ ( .D(n22754), .CK(clk), .Q(n19882), .QN(n28332) );
  DFF_X2 z_reg_2__7_ ( .D(n22775), .CK(clk), .Q(n20027), .QN(n28321) );
  DFF_X2 z_reg_2__6_ ( .D(n22783), .CK(clk), .Q(n20092), .QN(n28313) );
  DFF_X2 z_reg_2__4_ ( .D(n22799), .CK(clk), .Q(n20222), .QN(n28297) );
  DFF_X2 z_reg_63__14_ ( .D(n22947), .CK(clk), .Q(n19555), .QN(n28690) );
  DFF_X2 z_reg_63__7_ ( .D(n23017), .CK(clk), .Q(n20010), .QN(n28613) );
  DFF_X2 z_reg_63__6_ ( .D(n23027), .CK(clk), .Q(n20075), .QN(n28602) );
  DFF_X2 z_reg_63__5_ ( .D(n23037), .CK(clk), .Q(n20140), .QN(n28591) );
  DFF_X2 z_reg_63__1_ ( .D(n23077), .CK(clk), .Q(n20400), .QN(n28535) );
  DFF_X2 z_reg_63__13_ ( .D(n22957), .CK(clk), .Q(n19620), .QN(n28679) );
  DFF_X2 z_reg_63__12_ ( .D(n22967), .CK(clk), .Q(n19685), .QN(n28668) );
  DFF_X2 z_reg_63__11_ ( .D(n22977), .CK(clk), .Q(n19750), .QN(n28657) );
  DFF_X2 z_reg_63__10_ ( .D(n22987), .CK(clk), .Q(n19815), .QN(n28646) );
  DFF_X2 z_reg_63__9_ ( .D(n22997), .CK(clk), .Q(n19880), .QN(n28635) );
  DFF_X2 z_reg_63__8_ ( .D(n23007), .CK(clk), .Q(n19945), .QN(n28624) );
  DFF_X2 z_reg_63__4_ ( .D(n23047), .CK(clk), .Q(n20205), .QN(n28580) );
  DFF_X2 z_reg_63__3_ ( .D(n23057), .CK(clk), .Q(n20270), .QN(n28565) );
  DFF_X2 z_reg_63__2_ ( .D(n23067), .CK(clk), .Q(n20335), .QN(n28550) );
  DFF_X2 z_reg_63__0_ ( .D(n23087), .CK(clk), .Q(n20466), .QN(n28520) );
  DFF_X2 z_reg_53__12_ ( .D(n22607), .CK(clk), .Q(n19681), .QN(n28237) );
  DFF_X2 z_reg_53__9_ ( .D(n22631), .CK(clk), .Q(n19876), .QN(n28213) );
  DFF_X2 z_reg_53__8_ ( .D(n22639), .CK(clk), .Q(n19941), .QN(n28205) );
  DFF_X2 z_reg_53__7_ ( .D(n22647), .CK(clk), .Q(n20006), .QN(n28197) );
  DFF_X2 z_reg_53__6_ ( .D(n22655), .CK(clk), .Q(n20071), .QN(n28189) );
  DFF_X2 z_reg_53__5_ ( .D(n22663), .CK(clk), .Q(n20136), .QN(n28181) );
  DFF_X2 z_reg_53__4_ ( .D(n22671), .CK(clk), .Q(n20201), .QN(n28173) );
  DFF_X2 z_reg_53__3_ ( .D(n22679), .CK(clk), .Q(n20266), .QN(n28165) );
  DFF_X2 z_reg_53__2_ ( .D(n22687), .CK(clk), .Q(n20331), .QN(n28157) );
  DFF_X2 z_reg_53__1_ ( .D(n22695), .CK(clk), .Q(n20396), .QN(n28149) );
  DFF_X2 z_reg_53__0_ ( .D(n22703), .CK(clk), .Q(n20462), .QN(n28141) );
  DFF_X2 z_reg_42__14_ ( .D(n22941), .CK(clk), .Q(n19560), .QN(n28684) );
  DFF_X2 z_reg_42__13_ ( .D(n22951), .CK(clk), .Q(n19625), .QN(n28673) );
  DFF_X2 z_reg_42__12_ ( .D(n22961), .CK(clk), .Q(n19690), .QN(n28662) );
  DFF_X2 z_reg_42__11_ ( .D(n22971), .CK(clk), .Q(n19755), .QN(n28651) );
  DFF_X2 z_reg_42__10_ ( .D(n22981), .CK(clk), .Q(n19820), .QN(n28640) );
  DFF_X2 z_reg_42__9_ ( .D(n22991), .CK(clk), .Q(n19885), .QN(n28629) );
  DFF_X2 z_reg_42__8_ ( .D(n23001), .CK(clk), .Q(n19950), .QN(n28618) );
  DFF_X2 z_reg_42__7_ ( .D(n23011), .CK(clk), .Q(n20015), .QN(n28607) );
  DFF_X2 z_reg_42__6_ ( .D(n23021), .CK(clk), .Q(n20080), .QN(n28596) );
  DFF_X2 z_reg_42__5_ ( .D(n23031), .CK(clk), .Q(n20145), .QN(n28585) );
  DFF_X2 z_reg_42__4_ ( .D(n23041), .CK(clk), .Q(n20210), .QN(n28574) );
  DFF_X2 z_reg_42__3_ ( .D(n23051), .CK(clk), .Q(n20275), .QN(n28559) );
  DFF_X2 z_reg_42__2_ ( .D(n23061), .CK(clk), .Q(n20340), .QN(n28544) );
  DFF_X2 z_reg_42__1_ ( .D(n23071), .CK(clk), .Q(n20405), .QN(n28529) );
  DFF_X2 z_reg_42__0_ ( .D(n23081), .CK(clk), .Q(n20471), .QN(n28514) );
  DFF_X2 z_reg_34__8_ ( .D(n22763), .CK(clk), .Q(n19946), .QN(n28325) );
  DFF_X2 z_reg_34__7_ ( .D(n22771), .CK(clk), .Q(n20011), .QN(n28317) );
  DFF_X2 z_reg_34__6_ ( .D(n22779), .CK(clk), .Q(n20076), .QN(n28309) );
  DFF_X2 z_reg_34__5_ ( .D(n22787), .CK(clk), .Q(n20141), .QN(n28301) );
  DFF_X2 z_reg_34__4_ ( .D(n22795), .CK(clk), .Q(n20206), .QN(n28293) );
  DFF_X2 z_reg_34__3_ ( .D(n22803), .CK(clk), .Q(n20271), .QN(n28285) );
  DFF_X2 z_reg_34__2_ ( .D(n22811), .CK(clk), .Q(n20336), .QN(n28277) );
  DFF_X2 z_reg_34__1_ ( .D(n22819), .CK(clk), .Q(n20401), .QN(n28269) );
  DFF_X2 z_reg_34__0_ ( .D(n22827), .CK(clk), .Q(n20467), .QN(n28261) );
  DFF_X2 z_reg_24__14_ ( .D(n22841), .CK(clk), .Q(n19568), .QN(n28504) );
  DFF_X2 z_reg_24__13_ ( .D(n22847), .CK(clk), .Q(n19633), .QN(n28497) );
  DFF_X2 z_reg_24__12_ ( .D(n22853), .CK(clk), .Q(n19698), .QN(n28490) );
  DFF_X2 z_reg_24__11_ ( .D(n22859), .CK(clk), .Q(n19763), .QN(n28483) );
  DFF_X2 z_reg_24__10_ ( .D(n22865), .CK(clk), .Q(n19828), .QN(n28476) );
  DFF_X2 z_reg_24__9_ ( .D(n22871), .CK(clk), .Q(n19893), .QN(n28469) );
  DFF_X2 z_reg_24__8_ ( .D(n22877), .CK(clk), .Q(n19958), .QN(n28462) );
  DFF_X2 z_reg_24__7_ ( .D(n22883), .CK(clk), .Q(n20023), .QN(n28455) );
  DFF_X2 z_reg_24__6_ ( .D(n22889), .CK(clk), .Q(n20088), .QN(n28448) );
  DFF_X2 z_reg_24__5_ ( .D(n22895), .CK(clk), .Q(n20153), .QN(n28441) );
  DFF_X2 z_reg_24__4_ ( .D(n22901), .CK(clk), .Q(n20218), .QN(n28434) );
  DFF_X2 z_reg_24__3_ ( .D(n22907), .CK(clk), .Q(n20283), .QN(n28422) );
  DFF_X2 z_reg_24__2_ ( .D(n22913), .CK(clk), .Q(n20348), .QN(n28410) );
  DFF_X2 z_reg_24__1_ ( .D(n22919), .CK(clk), .Q(n20413), .QN(n28398) );
  DFF_X2 z_reg_24__0_ ( .D(n22925), .CK(clk), .Q(n20479), .QN(n28386) );
  DFF_X2 z_reg_16__8_ ( .D(n22635), .CK(clk), .Q(n19954), .QN(n28201) );
  DFF_X2 z_reg_16__7_ ( .D(n22643), .CK(clk), .Q(n20019), .QN(n28193) );
  DFF_X2 z_reg_16__6_ ( .D(n22651), .CK(clk), .Q(n20084), .QN(n28185) );
  DFF_X2 z_reg_16__5_ ( .D(n22659), .CK(clk), .Q(n20149), .QN(n28177) );
  DFF_X2 z_reg_16__4_ ( .D(n22667), .CK(clk), .Q(n20214), .QN(n28169) );
  DFF_X2 z_reg_16__3_ ( .D(n22675), .CK(clk), .Q(n20279), .QN(n28161) );
  DFF_X2 z_reg_16__2_ ( .D(n22683), .CK(clk), .Q(n20344), .QN(n28153) );
  DFF_X2 z_reg_16__1_ ( .D(n22691), .CK(clk), .Q(n20409), .QN(n28145) );
  DFF_X2 z_reg_16__0_ ( .D(n22699), .CK(clk), .Q(n20475), .QN(n28137) );
  DFF_X2 z_reg_48__14_ ( .D(n22590), .CK(clk), .Q(n19548), .QN(n28252) );
  DFF_X2 z_reg_48__13_ ( .D(n22598), .CK(clk), .Q(n19613), .QN(n28244) );
  DFF_X2 z_reg_48__12_ ( .D(n22606), .CK(clk), .Q(n19678), .QN(n28236) );
  DFF_X2 z_reg_48__11_ ( .D(n22614), .CK(clk), .Q(n19743), .QN(n28228) );
  DFF_X2 z_reg_48__10_ ( .D(n22622), .CK(clk), .Q(n19808), .QN(n28220) );
  DFF_X2 z_reg_48__9_ ( .D(n22630), .CK(clk), .Q(n19873), .QN(n28212) );
  DFF_X2 z_reg_2__14_ ( .D(n22719), .CK(clk), .Q(n19572), .QN(n28377) );
  DFF_X2 z_reg_2__13_ ( .D(n22727), .CK(clk), .Q(n19637), .QN(n28369) );
  DFF_X2 z_reg_2__12_ ( .D(n22735), .CK(clk), .Q(n19702), .QN(n28361) );
  DFF_X2 z_reg_2__11_ ( .D(n22743), .CK(clk), .Q(n19767), .QN(n28353) );
  DFF_X2 z_reg_2__10_ ( .D(n22751), .CK(clk), .Q(n19832), .QN(n28345) );
  DFF_X2 z_reg_2__9_ ( .D(n22759), .CK(clk), .Q(n19897), .QN(n28337) );
  DFF_X2 z_reg_53__14_ ( .D(n22591), .CK(clk), .Q(n19551), .QN(n28253) );
  DFF_X2 z_reg_53__13_ ( .D(n22599), .CK(clk), .Q(n19616), .QN(n28245) );
  DFF_X2 z_reg_53__11_ ( .D(n22615), .CK(clk), .Q(n19746), .QN(n28229) );
  DFF_X2 z_reg_53__10_ ( .D(n22623), .CK(clk), .Q(n19811), .QN(n28221) );
  DFF_X2 z_reg_16__14_ ( .D(n22587), .CK(clk), .Q(n19564), .QN(n28249) );
  DFF_X2 z_reg_16__13_ ( .D(n22595), .CK(clk), .Q(n19629), .QN(n28241) );
  DFF_X2 z_reg_16__12_ ( .D(n22603), .CK(clk), .Q(n19694), .QN(n28233) );
  DFF_X2 z_reg_16__11_ ( .D(n22611), .CK(clk), .Q(n19759), .QN(n28225) );
  DFF_X2 z_reg_16__10_ ( .D(n22619), .CK(clk), .Q(n19824), .QN(n28217) );
  DFF_X2 z_reg_16__9_ ( .D(n22627), .CK(clk), .Q(n19889), .QN(n28209) );
  DFF_X2 z_reg_34__14_ ( .D(n22715), .CK(clk), .Q(n19556), .QN(n28373) );
  DFF_X2 z_reg_34__13_ ( .D(n22723), .CK(clk), .Q(n19621), .QN(n28365) );
  DFF_X2 z_reg_34__12_ ( .D(n22731), .CK(clk), .Q(n19686), .QN(n28357) );
  DFF_X2 z_reg_34__11_ ( .D(n22739), .CK(clk), .Q(n19751), .QN(n28349) );
  DFF_X2 z_reg_34__10_ ( .D(n22747), .CK(clk), .Q(n19816), .QN(n28341) );
  DFF_X2 z_reg_34__9_ ( .D(n22755), .CK(clk), .Q(n19881), .QN(n28333) );
  DFF_X2 z_reg_47__14_ ( .D(n22938), .CK(clk), .QN(n28681) );
  DFF_X2 z_reg_47__13_ ( .D(n22948), .CK(clk), .QN(n28670) );
  DFF_X2 z_reg_47__12_ ( .D(n22958), .CK(clk), .QN(n28659) );
  DFF_X2 z_reg_47__11_ ( .D(n22968), .CK(clk), .QN(n28648) );
  DFF_X2 z_reg_47__10_ ( .D(n22978), .CK(clk), .QN(n28637) );
  DFF_X2 z_reg_47__9_ ( .D(n22988), .CK(clk), .QN(n28626) );
  DFF_X2 z_reg_47__8_ ( .D(n22998), .CK(clk), .QN(n28615) );
  DFF_X2 z_reg_47__7_ ( .D(n23008), .CK(clk), .QN(n28604) );
  DFF_X2 z_reg_47__6_ ( .D(n23018), .CK(clk), .QN(n28593) );
  DFF_X2 z_reg_47__5_ ( .D(n23028), .CK(clk), .QN(n28582) );
  DFF_X2 z_reg_47__4_ ( .D(n23038), .CK(clk), .QN(n28571) );
  DFF_X2 z_reg_47__3_ ( .D(n23048), .CK(clk), .QN(n28556) );
  DFF_X2 z_reg_47__2_ ( .D(n23058), .CK(clk), .QN(n28541) );
  DFF_X2 z_reg_47__1_ ( .D(n23068), .CK(clk), .QN(n28526) );
  DFF_X2 z_reg_47__0_ ( .D(n23078), .CK(clk), .QN(n28511) );
  DFF_X2 z_reg_39__8_ ( .D(n22760), .CK(clk), .QN(n28322) );
  DFF_X2 z_reg_39__7_ ( .D(n22768), .CK(clk), .QN(n28314) );
  DFF_X2 z_reg_39__6_ ( .D(n22776), .CK(clk), .QN(n28306) );
  DFF_X2 z_reg_39__5_ ( .D(n22784), .CK(clk), .QN(n28298) );
  DFF_X2 z_reg_39__4_ ( .D(n22792), .CK(clk), .QN(n28290) );
  DFF_X2 z_reg_39__3_ ( .D(n22800), .CK(clk), .QN(n28282) );
  DFF_X2 z_reg_39__2_ ( .D(n22808), .CK(clk), .QN(n28274) );
  DFF_X2 z_reg_39__1_ ( .D(n22816), .CK(clk), .QN(n28266) );
  DFF_X2 z_reg_39__0_ ( .D(n22824), .CK(clk), .QN(n28258) );
  DFF_X2 z_reg_29__14_ ( .D(n22838), .CK(clk), .QN(n28501) );
  DFF_X2 z_reg_29__13_ ( .D(n22844), .CK(clk), .QN(n28494) );
  DFF_X2 z_reg_29__12_ ( .D(n22850), .CK(clk), .QN(n28487) );
  DFF_X2 z_reg_29__11_ ( .D(n22856), .CK(clk), .QN(n28480) );
  DFF_X2 z_reg_29__10_ ( .D(n22862), .CK(clk), .QN(n28473) );
  DFF_X2 z_reg_29__9_ ( .D(n22868), .CK(clk), .QN(n28466) );
  DFF_X2 z_reg_29__8_ ( .D(n22874), .CK(clk), .QN(n28459) );
  DFF_X2 z_reg_29__7_ ( .D(n22880), .CK(clk), .QN(n28452) );
  DFF_X2 z_reg_29__6_ ( .D(n22886), .CK(clk), .QN(n28445) );
  DFF_X2 z_reg_29__5_ ( .D(n22892), .CK(clk), .QN(n28438) );
  DFF_X2 z_reg_29__4_ ( .D(n22898), .CK(clk), .QN(n28431) );
  DFF_X2 z_reg_29__3_ ( .D(n22904), .CK(clk), .QN(n28419) );
  DFF_X2 z_reg_29__2_ ( .D(n22910), .CK(clk), .QN(n28407) );
  DFF_X2 z_reg_29__1_ ( .D(n22916), .CK(clk), .QN(n28395) );
  DFF_X2 z_reg_29__0_ ( .D(n22922), .CK(clk), .QN(n28383) );
  DFF_X2 z_reg_21__8_ ( .D(n22632), .CK(clk), .QN(n28198) );
  DFF_X2 z_reg_21__7_ ( .D(n22640), .CK(clk), .QN(n28190) );
  DFF_X2 z_reg_21__6_ ( .D(n22648), .CK(clk), .QN(n28182) );
  DFF_X2 z_reg_21__5_ ( .D(n22656), .CK(clk), .QN(n28174) );
  DFF_X2 z_reg_21__4_ ( .D(n22664), .CK(clk), .QN(n28166) );
  DFF_X2 z_reg_21__3_ ( .D(n22672), .CK(clk), .QN(n28158) );
  DFF_X2 z_reg_21__2_ ( .D(n22680), .CK(clk), .QN(n28150) );
  DFF_X2 z_reg_21__1_ ( .D(n22688), .CK(clk), .QN(n28142) );
  DFF_X2 z_reg_21__0_ ( .D(n22696), .CK(clk), .QN(n28134) );
  DFF_X2 z_reg_15__14_ ( .D(n22945), .CK(clk), .Q(n19579), .QN(n28688) );
  DFF_X2 z_reg_15__13_ ( .D(n22955), .CK(clk), .Q(n19644), .QN(n28677) );
  DFF_X2 z_reg_15__12_ ( .D(n22965), .CK(clk), .Q(n19709), .QN(n28666) );
  DFF_X2 z_reg_15__11_ ( .D(n22975), .CK(clk), .Q(n19774), .QN(n28655) );
  DFF_X2 z_reg_15__10_ ( .D(n22985), .CK(clk), .Q(n19839), .QN(n28644) );
  DFF_X2 z_reg_15__9_ ( .D(n22995), .CK(clk), .Q(n19904), .QN(n28633) );
  DFF_X2 z_reg_15__8_ ( .D(n23005), .CK(clk), .Q(n19969), .QN(n28622) );
  DFF_X2 z_reg_15__7_ ( .D(n23015), .CK(clk), .Q(n20034), .QN(n28611) );
  DFF_X2 z_reg_15__6_ ( .D(n23025), .CK(clk), .Q(n20099), .QN(n28600) );
  DFF_X2 z_reg_15__5_ ( .D(n23035), .CK(clk), .Q(n20164), .QN(n28589) );
  DFF_X2 z_reg_15__4_ ( .D(n23045), .CK(clk), .Q(n20229), .QN(n28578) );
  DFF_X2 z_reg_15__3_ ( .D(n23055), .CK(clk), .Q(n20294), .QN(n28563) );
  DFF_X2 z_reg_15__2_ ( .D(n23065), .CK(clk), .Q(n20359), .QN(n28548) );
  DFF_X2 z_reg_15__1_ ( .D(n23075), .CK(clk), .Q(n20424), .QN(n28533) );
  DFF_X2 z_reg_15__0_ ( .D(n23085), .CK(clk), .Q(n20490), .QN(n28518) );
  DFF_X2 z_reg_7__8_ ( .D(n22766), .CK(clk), .QN(n28328) );
  DFF_X2 z_reg_7__7_ ( .D(n22774), .CK(clk), .QN(n28320) );
  DFF_X2 z_reg_7__6_ ( .D(n22782), .CK(clk), .QN(n28312) );
  DFF_X2 z_reg_7__5_ ( .D(n22790), .CK(clk), .QN(n28304) );
  DFF_X2 z_reg_7__4_ ( .D(n22798), .CK(clk), .QN(n28296) );
  DFF_X2 z_reg_7__3_ ( .D(n22806), .CK(clk), .QN(n28288) );
  DFF_X2 z_reg_7__2_ ( .D(n22814), .CK(clk), .QN(n28280) );
  DFF_X2 z_reg_7__1_ ( .D(n22822), .CK(clk), .QN(n28272) );
  DFF_X2 z_reg_7__0_ ( .D(n22830), .CK(clk), .QN(n28264) );
  DFF_X2 z_reg_39__14_ ( .D(n22712), .CK(clk), .QN(n28370) );
  DFF_X2 z_reg_39__13_ ( .D(n22720), .CK(clk), .QN(n28362) );
  DFF_X2 z_reg_39__12_ ( .D(n22728), .CK(clk), .QN(n28354) );
  DFF_X2 z_reg_39__11_ ( .D(n22736), .CK(clk), .QN(n28346) );
  DFF_X2 z_reg_39__10_ ( .D(n22744), .CK(clk), .QN(n28338) );
  DFF_X2 z_reg_39__9_ ( .D(n22752), .CK(clk), .QN(n28330) );
  DFF_X2 z_reg_21__14_ ( .D(n22584), .CK(clk), .QN(n28246) );
  DFF_X2 z_reg_21__13_ ( .D(n22592), .CK(clk), .QN(n28238) );
  DFF_X2 z_reg_21__12_ ( .D(n22600), .CK(clk), .QN(n28230) );
  DFF_X2 z_reg_21__11_ ( .D(n22608), .CK(clk), .QN(n28222) );
  DFF_X2 z_reg_21__10_ ( .D(n22616), .CK(clk), .QN(n28214) );
  DFF_X2 z_reg_21__9_ ( .D(n22624), .CK(clk), .QN(n28206) );
  DFF_X2 z_reg_7__14_ ( .D(n22718), .CK(clk), .QN(n28376) );
  DFF_X2 z_reg_7__13_ ( .D(n22726), .CK(clk), .QN(n28368) );
  DFF_X2 z_reg_7__12_ ( .D(n22734), .CK(clk), .QN(n28360) );
  DFF_X2 z_reg_7__11_ ( .D(n22742), .CK(clk), .QN(n28352) );
  DFF_X2 z_reg_7__10_ ( .D(n22750), .CK(clk), .QN(n28344) );
  DFF_X2 z_reg_7__9_ ( .D(n22758), .CK(clk), .QN(n28336) );
  DFF_X2 output_store_reg_6__15_ ( .D(n25262), .CK(clk), .Q(n26166), .QN(
        n28817) );
  DFF_X2 output_store_reg_4__15_ ( .D(n24898), .CK(clk), .Q(n19355) );
  DFF_X2 output_store_reg_3__15_ ( .D(n24897), .CK(clk), .Q(n19356) );
  DFF_X2 output_store_reg_2__15_ ( .D(n25260), .CK(clk), .Q(n26164), .QN(
        n28819) );
  DFF_X2 output_store_reg_1__15_ ( .D(n25259), .CK(clk), .Q(n26163), .QN(
        n28820) );
  DFF_X2 output_store_reg_0__15_ ( .D(n25258), .CK(clk), .Q(n26162), .QN(
        n28821) );
  DFF_X2 output_store_reg_5__14_ ( .D(n22458), .CK(clk), .QN(n28811) );
  DFF_X2 output_store_reg_5__13_ ( .D(n22466), .CK(clk), .QN(n28803) );
  DFF_X2 output_store_reg_5__12_ ( .D(n22474), .CK(clk), .QN(n28795) );
  DFF_X2 output_store_reg_5__11_ ( .D(n22482), .CK(clk), .QN(n28787) );
  DFF_X2 output_store_reg_5__10_ ( .D(n22490), .CK(clk), .QN(n28779) );
  DFF_X2 output_store_reg_5__9_ ( .D(n22498), .CK(clk), .QN(n28771) );
  DFF_X2 output_store_reg_5__8_ ( .D(n22506), .CK(clk), .QN(n28763) );
  DFF_X2 output_store_reg_5__4_ ( .D(n22538), .CK(clk), .QN(n28731) );
  DFF_X2 output_store_reg_5__3_ ( .D(n22546), .CK(clk), .QN(n28723) );
  DFF_X2 output_store_reg_5__2_ ( .D(n22554), .CK(clk), .QN(n28715) );
  DFF_X2 output_store_reg_5__0_ ( .D(n22570), .CK(clk), .QN(n28699) );
  DFF_X2 output_store_reg_5__7_ ( .D(n22514), .CK(clk), .QN(n28755) );
  DFF_X2 output_store_reg_5__6_ ( .D(n22522), .CK(clk), .QN(n28747) );
  DFF_X2 output_store_reg_5__5_ ( .D(n22530), .CK(clk), .QN(n28739) );
  DFF_X2 output_store_reg_5__1_ ( .D(n22562), .CK(clk), .QN(n28707) );
  DFF_X2 count_out_reg_0_ ( .D(n23433), .CK(clk), .Q(n19348), .QN(n26129) );
  DFF_X2 output_store_reg_6__14_ ( .D(n22457), .CK(clk), .QN(n28810) );
  DFF_X2 output_store_reg_6__13_ ( .D(n22465), .CK(clk), .QN(n28802) );
  DFF_X2 output_store_reg_6__12_ ( .D(n22473), .CK(clk), .QN(n28794) );
  DFF_X2 output_store_reg_6__11_ ( .D(n22481), .CK(clk), .QN(n28786) );
  DFF_X2 output_store_reg_6__10_ ( .D(n22489), .CK(clk), .QN(n28778) );
  DFF_X2 output_store_reg_6__9_ ( .D(n22497), .CK(clk), .QN(n28770) );
  DFF_X2 output_store_reg_6__8_ ( .D(n22505), .CK(clk), .QN(n28762) );
  DFF_X2 output_store_reg_6__7_ ( .D(n22513), .CK(clk), .QN(n28754) );
  DFF_X2 output_store_reg_6__6_ ( .D(n22521), .CK(clk), .QN(n28746) );
  DFF_X2 output_store_reg_6__5_ ( .D(n22529), .CK(clk), .QN(n28738) );
  DFF_X2 output_store_reg_6__4_ ( .D(n22537), .CK(clk), .QN(n28730) );
  DFF_X2 output_store_reg_6__3_ ( .D(n22545), .CK(clk), .QN(n28722) );
  DFF_X2 output_store_reg_6__2_ ( .D(n22553), .CK(clk), .QN(n28714) );
  DFF_X2 output_store_reg_6__1_ ( .D(n22561), .CK(clk), .QN(n28706) );
  DFF_X2 output_store_reg_6__0_ ( .D(n22569), .CK(clk), .QN(n28698) );
  DFF_X2 output_store_reg_7__14_ ( .D(n22456), .CK(clk), .Q(n19360), .QN(
        n28809) );
  DFF_X2 output_store_reg_7__13_ ( .D(n22464), .CK(clk), .Q(n19368), .QN(
        n28801) );
  DFF_X2 output_store_reg_7__12_ ( .D(n22472), .CK(clk), .Q(n19376), .QN(
        n28793) );
  DFF_X2 output_store_reg_7__11_ ( .D(n22480), .CK(clk), .Q(n19384), .QN(
        n28785) );
  DFF_X2 output_store_reg_7__10_ ( .D(n22488), .CK(clk), .Q(n19392), .QN(
        n28777) );
  DFF_X2 output_store_reg_7__9_ ( .D(n22496), .CK(clk), .Q(n19400), .QN(n28769) );
  DFF_X2 output_store_reg_7__8_ ( .D(n22504), .CK(clk), .Q(n19408), .QN(n28761) );
  DFF_X2 output_store_reg_7__7_ ( .D(n22512), .CK(clk), .Q(n19416), .QN(n28753) );
  DFF_X2 output_store_reg_7__6_ ( .D(n22520), .CK(clk), .Q(n19424), .QN(n28745) );
  DFF_X2 output_store_reg_7__5_ ( .D(n22528), .CK(clk), .Q(n19432), .QN(n28737) );
  DFF_X2 output_store_reg_7__4_ ( .D(n22536), .CK(clk), .Q(n19440), .QN(n28729) );
  DFF_X2 output_store_reg_7__3_ ( .D(n22544), .CK(clk), .Q(n19448), .QN(n28721) );
  DFF_X2 output_store_reg_7__2_ ( .D(n22552), .CK(clk), .Q(n19456), .QN(n28713) );
  DFF_X2 output_store_reg_7__1_ ( .D(n22560), .CK(clk), .Q(n19464), .QN(n28705) );
  DFF_X2 output_store_reg_7__0_ ( .D(n22568), .CK(clk), .Q(n19472), .QN(n28697) );
  DFF_X2 output_store_reg_4__14_ ( .D(n22459), .CK(clk), .Q(n19363), .QN(
        n28812) );
  DFF_X2 output_store_reg_4__13_ ( .D(n22467), .CK(clk), .Q(n19371), .QN(
        n28804) );
  DFF_X2 output_store_reg_4__12_ ( .D(n22475), .CK(clk), .Q(n19379), .QN(
        n28796) );
  DFF_X2 output_store_reg_4__11_ ( .D(n22483), .CK(clk), .Q(n19387), .QN(
        n28788) );
  DFF_X2 output_store_reg_4__10_ ( .D(n22491), .CK(clk), .Q(n19395), .QN(
        n28780) );
  DFF_X2 output_store_reg_4__9_ ( .D(n22499), .CK(clk), .Q(n19403), .QN(n28772) );
  DFF_X2 output_store_reg_4__8_ ( .D(n22507), .CK(clk), .Q(n19411), .QN(n28764) );
  DFF_X2 output_store_reg_4__4_ ( .D(n22539), .CK(clk), .Q(n19443), .QN(n28732) );
  DFF_X2 output_store_reg_4__3_ ( .D(n22547), .CK(clk), .Q(n19451), .QN(n28724) );
  DFF_X2 output_store_reg_4__2_ ( .D(n22555), .CK(clk), .Q(n19459), .QN(n28716) );
  DFF_X2 output_store_reg_4__0_ ( .D(n22571), .CK(clk), .Q(n19475), .QN(n28700) );
  DFF_X2 output_store_reg_4__7_ ( .D(n22515), .CK(clk), .Q(n19419), .QN(n28756) );
  DFF_X2 output_store_reg_4__6_ ( .D(n22523), .CK(clk), .Q(n19427), .QN(n28748) );
  DFF_X2 output_store_reg_4__5_ ( .D(n22531), .CK(clk), .Q(n19435), .QN(n28740) );
  DFF_X2 output_store_reg_4__1_ ( .D(n22563), .CK(clk), .Q(n19467), .QN(n28708) );
  DFF_X2 output_store_reg_7__15_ ( .D(n24893), .CK(clk), .Q(n19352) );
  DFF_X2 output_store_reg_3__14_ ( .D(n22460), .CK(clk), .Q(n19364), .QN(
        n28813) );
  DFF_X2 output_store_reg_3__13_ ( .D(n22468), .CK(clk), .Q(n19372), .QN(
        n28805) );
  DFF_X2 output_store_reg_3__12_ ( .D(n22476), .CK(clk), .Q(n19380), .QN(
        n28797) );
  DFF_X2 output_store_reg_3__11_ ( .D(n22484), .CK(clk), .Q(n19388), .QN(
        n28789) );
  DFF_X2 output_store_reg_3__10_ ( .D(n22492), .CK(clk), .Q(n19396), .QN(
        n28781) );
  DFF_X2 output_store_reg_3__9_ ( .D(n22500), .CK(clk), .Q(n19404), .QN(n28773) );
  DFF_X2 output_store_reg_3__8_ ( .D(n22508), .CK(clk), .Q(n19412), .QN(n28765) );
  DFF_X2 output_store_reg_3__4_ ( .D(n22540), .CK(clk), .Q(n19444), .QN(n28733) );
  DFF_X2 output_store_reg_3__3_ ( .D(n22548), .CK(clk), .Q(n19452), .QN(n28725) );
  DFF_X2 output_store_reg_3__2_ ( .D(n22556), .CK(clk), .Q(n19460), .QN(n28717) );
  DFF_X2 output_store_reg_3__0_ ( .D(n22572), .CK(clk), .Q(n19476), .QN(n28701) );
  DFF_X2 output_store_reg_2__14_ ( .D(n22461), .CK(clk), .QN(n28814) );
  DFF_X2 output_store_reg_2__13_ ( .D(n22469), .CK(clk), .QN(n28806) );
  DFF_X2 output_store_reg_2__12_ ( .D(n22477), .CK(clk), .QN(n28798) );
  DFF_X2 output_store_reg_2__11_ ( .D(n22485), .CK(clk), .QN(n28790) );
  DFF_X2 output_store_reg_2__10_ ( .D(n22493), .CK(clk), .QN(n28782) );
  DFF_X2 output_store_reg_2__9_ ( .D(n22501), .CK(clk), .QN(n28774) );
  DFF_X2 output_store_reg_2__8_ ( .D(n22509), .CK(clk), .QN(n28766) );
  DFF_X2 output_store_reg_2__4_ ( .D(n22541), .CK(clk), .QN(n28734) );
  DFF_X2 output_store_reg_2__3_ ( .D(n22549), .CK(clk), .QN(n28726) );
  DFF_X2 output_store_reg_2__2_ ( .D(n22557), .CK(clk), .QN(n28718) );
  DFF_X2 output_store_reg_2__0_ ( .D(n22573), .CK(clk), .QN(n28702) );
  DFF_X2 output_store_reg_1__14_ ( .D(n22462), .CK(clk), .QN(n28815) );
  DFF_X2 output_store_reg_1__13_ ( .D(n22470), .CK(clk), .QN(n28807) );
  DFF_X2 output_store_reg_1__12_ ( .D(n22478), .CK(clk), .QN(n28799) );
  DFF_X2 output_store_reg_1__11_ ( .D(n22486), .CK(clk), .QN(n28791) );
  DFF_X2 output_store_reg_1__10_ ( .D(n22494), .CK(clk), .QN(n28783) );
  DFF_X2 output_store_reg_1__9_ ( .D(n22502), .CK(clk), .QN(n28775) );
  DFF_X2 output_store_reg_1__8_ ( .D(n22510), .CK(clk), .QN(n28767) );
  DFF_X2 output_store_reg_1__4_ ( .D(n22542), .CK(clk), .QN(n28735) );
  DFF_X2 output_store_reg_1__3_ ( .D(n22550), .CK(clk), .QN(n28727) );
  DFF_X2 output_store_reg_1__2_ ( .D(n22558), .CK(clk), .QN(n28719) );
  DFF_X2 output_store_reg_1__0_ ( .D(n22574), .CK(clk), .QN(n28703) );
  DFF_X2 output_store_reg_0__14_ ( .D(n22463), .CK(clk), .QN(n28816) );
  DFF_X2 output_store_reg_0__13_ ( .D(n22471), .CK(clk), .QN(n28808) );
  DFF_X2 output_store_reg_0__12_ ( .D(n22479), .CK(clk), .QN(n28800) );
  DFF_X2 output_store_reg_0__11_ ( .D(n22487), .CK(clk), .QN(n28792) );
  DFF_X2 output_store_reg_0__10_ ( .D(n22495), .CK(clk), .QN(n28784) );
  DFF_X2 output_store_reg_0__9_ ( .D(n22503), .CK(clk), .QN(n28776) );
  DFF_X2 output_store_reg_0__8_ ( .D(n22511), .CK(clk), .QN(n28768) );
  DFF_X2 output_store_reg_0__4_ ( .D(n22543), .CK(clk), .QN(n28736) );
  DFF_X2 output_store_reg_0__3_ ( .D(n22551), .CK(clk), .QN(n28728) );
  DFF_X2 output_store_reg_0__2_ ( .D(n22559), .CK(clk), .QN(n28720) );
  DFF_X2 output_store_reg_0__0_ ( .D(n22575), .CK(clk), .QN(n28704) );
  DFF_X2 output_store_reg_3__7_ ( .D(n22516), .CK(clk), .Q(n19420), .QN(n28757) );
  DFF_X2 output_store_reg_3__6_ ( .D(n22524), .CK(clk), .Q(n19428), .QN(n28749) );
  DFF_X2 output_store_reg_3__5_ ( .D(n22532), .CK(clk), .Q(n19436), .QN(n28741) );
  DFF_X2 output_store_reg_3__1_ ( .D(n22564), .CK(clk), .Q(n19468), .QN(n28709) );
  DFF_X2 output_store_reg_2__7_ ( .D(n22517), .CK(clk), .QN(n28758) );
  DFF_X2 output_store_reg_2__6_ ( .D(n22525), .CK(clk), .QN(n28750) );
  DFF_X2 output_store_reg_2__5_ ( .D(n22533), .CK(clk), .QN(n28742) );
  DFF_X2 output_store_reg_2__1_ ( .D(n22565), .CK(clk), .QN(n28710) );
  DFF_X2 output_store_reg_1__7_ ( .D(n22518), .CK(clk), .QN(n28759) );
  DFF_X2 output_store_reg_1__6_ ( .D(n22526), .CK(clk), .QN(n28751) );
  DFF_X2 output_store_reg_1__5_ ( .D(n22534), .CK(clk), .QN(n28743) );
  DFF_X2 output_store_reg_1__1_ ( .D(n22566), .CK(clk), .QN(n28711) );
  DFF_X2 output_store_reg_0__7_ ( .D(n22519), .CK(clk), .QN(n28760) );
  DFF_X2 output_store_reg_0__6_ ( .D(n22527), .CK(clk), .QN(n28752) );
  DFF_X2 output_store_reg_0__5_ ( .D(n22535), .CK(clk), .QN(n28744) );
  DFF_X2 output_store_reg_0__1_ ( .D(n22567), .CK(clk), .QN(n28712) );
  DFF_X2 count_store_reg_3_ ( .D(n24819), .CK(clk), .Q(n19349), .QN(n28822) );
  DFF_X2 bitselect2_reg_3_ ( .D(n23447), .CK(clk), .Q(n18743), .QN(n26136) );
  DFF_X2 dut__dom__data_reg_15_ ( .D(n22446), .CK(clk), .Q(dut__dom__data[15])
         );
  DFF_X2 dut__dom__data_reg_14_ ( .D(n22445), .CK(clk), .Q(dut__dom__data[14])
         );
  DFF_X2 dut__dom__data_reg_13_ ( .D(n22444), .CK(clk), .Q(dut__dom__data[13])
         );
  DFF_X2 dut__dom__data_reg_12_ ( .D(n22443), .CK(clk), .Q(dut__dom__data[12])
         );
  DFF_X2 dut__dom__data_reg_11_ ( .D(n22442), .CK(clk), .Q(dut__dom__data[11])
         );
  DFF_X2 dut__dom__data_reg_10_ ( .D(n22441), .CK(clk), .Q(dut__dom__data[10])
         );
  DFF_X2 dut__dom__data_reg_9_ ( .D(n22440), .CK(clk), .Q(dut__dom__data[9])
         );
  DFF_X2 dut__dom__data_reg_8_ ( .D(n22439), .CK(clk), .Q(dut__dom__data[8])
         );
  DFF_X2 dut__dom__data_reg_7_ ( .D(n22438), .CK(clk), .Q(dut__dom__data[7])
         );
  DFF_X2 dut__dom__data_reg_6_ ( .D(n22437), .CK(clk), .Q(dut__dom__data[6])
         );
  DFF_X2 dut__dom__data_reg_5_ ( .D(n22436), .CK(clk), .Q(dut__dom__data[5])
         );
  DFF_X2 dut__dom__data_reg_4_ ( .D(n22435), .CK(clk), .Q(dut__dom__data[4])
         );
  DFF_X2 dut__dom__data_reg_3_ ( .D(n22434), .CK(clk), .Q(dut__dom__data[3])
         );
  DFF_X2 dut__dom__data_reg_2_ ( .D(n22433), .CK(clk), .Q(dut__dom__data[2])
         );
  DFF_X2 dut__dom__data_reg_1_ ( .D(n22432), .CK(clk), .Q(dut__dom__data[1])
         );
  DFF_X2 dut__dom__data_reg_0_ ( .D(n22431), .CK(clk), .Q(dut__dom__data[0])
         );
  DFF_X2 avector30_reg_0__15_ ( .D(n24809), .CK(clk), .Q(n16394), .QN(n27542)
         );
  DFF_X2 avector30_reg_0__14_ ( .D(n24808), .CK(clk), .Q(n16431), .QN(n27541)
         );
  DFF_X2 avector30_reg_0__13_ ( .D(n24807), .CK(clk), .Q(n16468), .QN(n27540)
         );
  DFF_X2 avector30_reg_0__12_ ( .D(n24806), .CK(clk), .Q(n16505), .QN(n27539)
         );
  DFF_X2 avector30_reg_0__11_ ( .D(n24805), .CK(clk), .Q(n16542), .QN(n27538)
         );
  DFF_X2 avector30_reg_0__10_ ( .D(n24804), .CK(clk), .Q(n16579), .QN(n27537)
         );
  DFF_X2 avector30_reg_0__9_ ( .D(n24803), .CK(clk), .Q(n16616), .QN(n27536)
         );
  DFF_X2 avector30_reg_0__8_ ( .D(n24802), .CK(clk), .Q(n16653), .QN(n27535)
         );
  DFF_X2 avector30_reg_0__7_ ( .D(n24801), .CK(clk), .Q(n16690), .QN(n27534)
         );
  DFF_X2 avector30_reg_0__6_ ( .D(n24800), .CK(clk), .Q(n16727), .QN(n27533)
         );
  DFF_X2 avector30_reg_0__5_ ( .D(n24799), .CK(clk), .Q(n16764), .QN(n27532)
         );
  DFF_X2 avector30_reg_0__4_ ( .D(n24798), .CK(clk), .Q(n16801), .QN(n27531)
         );
  DFF_X2 avector30_reg_0__3_ ( .D(n24797), .CK(clk), .Q(n16838), .QN(n27530)
         );
  DFF_X2 avector30_reg_0__2_ ( .D(n24796), .CK(clk), .Q(n16875), .QN(n27529)
         );
  DFF_X2 avector30_reg_0__1_ ( .D(n24795), .CK(clk), .Q(n16912), .QN(n27528)
         );
  DFF_X2 avector30_reg_0__0_ ( .D(n24794), .CK(clk), .Q(n16949), .QN(n27527)
         );
  DFF_X2 avector32_reg_8__15_ ( .D(n24099), .CK(clk), .QN(n26550) );
  DFF_X2 avector32_reg_8__14_ ( .D(n24098), .CK(clk), .QN(n26549) );
  DFF_X2 avector32_reg_8__13_ ( .D(n24097), .CK(clk), .QN(n26548) );
  DFF_X2 avector32_reg_8__12_ ( .D(n24096), .CK(clk), .QN(n26547) );
  DFF_X2 avector32_reg_8__11_ ( .D(n24095), .CK(clk), .QN(n26546) );
  DFF_X2 avector32_reg_8__10_ ( .D(n24094), .CK(clk), .QN(n26545) );
  DFF_X2 avector32_reg_8__9_ ( .D(n24093), .CK(clk), .QN(n26544) );
  DFF_X2 avector32_reg_8__8_ ( .D(n24092), .CK(clk), .QN(n26543) );
  DFF_X2 avector32_reg_8__7_ ( .D(n24091), .CK(clk), .QN(n26542) );
  DFF_X2 avector32_reg_8__6_ ( .D(n24090), .CK(clk), .QN(n26541) );
  DFF_X2 avector32_reg_8__5_ ( .D(n24089), .CK(clk), .QN(n26540) );
  DFF_X2 avector32_reg_8__4_ ( .D(n24088), .CK(clk), .QN(n26539) );
  DFF_X2 avector32_reg_8__3_ ( .D(n24087), .CK(clk), .QN(n26538) );
  DFF_X2 avector32_reg_8__2_ ( .D(n24086), .CK(clk), .QN(n26537) );
  DFF_X2 avector32_reg_8__1_ ( .D(n24085), .CK(clk), .QN(n26536) );
  DFF_X2 avector32_reg_8__0_ ( .D(n24084), .CK(clk), .QN(n26535) );
  DFF_X2 avector31_reg_8__15_ ( .D(n24419), .CK(clk), .QN(n26646) );
  DFF_X2 avector31_reg_8__14_ ( .D(n24418), .CK(clk), .QN(n26645) );
  DFF_X2 avector31_reg_8__13_ ( .D(n24417), .CK(clk), .QN(n26644) );
  DFF_X2 avector31_reg_8__12_ ( .D(n24416), .CK(clk), .QN(n26643) );
  DFF_X2 avector31_reg_8__11_ ( .D(n24415), .CK(clk), .QN(n26642) );
  DFF_X2 avector31_reg_8__10_ ( .D(n24414), .CK(clk), .QN(n26641) );
  DFF_X2 avector31_reg_8__9_ ( .D(n24413), .CK(clk), .QN(n26640) );
  DFF_X2 avector31_reg_8__8_ ( .D(n24412), .CK(clk), .QN(n26639) );
  DFF_X2 avector31_reg_8__7_ ( .D(n24411), .CK(clk), .QN(n26638) );
  DFF_X2 avector31_reg_8__6_ ( .D(n24410), .CK(clk), .QN(n26637) );
  DFF_X2 avector31_reg_8__5_ ( .D(n24409), .CK(clk), .QN(n26636) );
  DFF_X2 avector31_reg_8__4_ ( .D(n24408), .CK(clk), .QN(n26635) );
  DFF_X2 avector31_reg_8__3_ ( .D(n24407), .CK(clk), .QN(n26634) );
  DFF_X2 avector31_reg_8__2_ ( .D(n24406), .CK(clk), .QN(n26633) );
  DFF_X2 avector31_reg_8__1_ ( .D(n24405), .CK(clk), .QN(n26632) );
  DFF_X2 avector31_reg_8__0_ ( .D(n24404), .CK(clk), .QN(n26631) );
  DFF_X2 avector30_reg_8__15_ ( .D(n24745), .CK(clk), .Q(n16398), .QN(n26614)
         );
  DFF_X2 avector30_reg_8__14_ ( .D(n24744), .CK(clk), .Q(n16435), .QN(n26613)
         );
  DFF_X2 avector30_reg_8__13_ ( .D(n24743), .CK(clk), .Q(n16472), .QN(n26612)
         );
  DFF_X2 avector30_reg_8__12_ ( .D(n24742), .CK(clk), .Q(n16509), .QN(n26611)
         );
  DFF_X2 avector30_reg_8__11_ ( .D(n24741), .CK(clk), .Q(n16546), .QN(n26610)
         );
  DFF_X2 avector30_reg_8__10_ ( .D(n24740), .CK(clk), .Q(n16583), .QN(n26609)
         );
  DFF_X2 avector30_reg_8__9_ ( .D(n24739), .CK(clk), .Q(n16620), .QN(n26608)
         );
  DFF_X2 avector30_reg_8__8_ ( .D(n24738), .CK(clk), .Q(n16657), .QN(n26607)
         );
  DFF_X2 avector30_reg_8__7_ ( .D(n24737), .CK(clk), .Q(n16694), .QN(n26606)
         );
  DFF_X2 avector30_reg_8__6_ ( .D(n24736), .CK(clk), .Q(n16731), .QN(n26605)
         );
  DFF_X2 avector30_reg_8__5_ ( .D(n24735), .CK(clk), .Q(n16768), .QN(n26604)
         );
  DFF_X2 avector30_reg_8__4_ ( .D(n24734), .CK(clk), .Q(n16805), .QN(n26603)
         );
  DFF_X2 avector30_reg_8__3_ ( .D(n24733), .CK(clk), .Q(n16842), .QN(n26602)
         );
  DFF_X2 avector30_reg_8__2_ ( .D(n24732), .CK(clk), .Q(n16879), .QN(n26601)
         );
  DFF_X2 avector30_reg_8__1_ ( .D(n24731), .CK(clk), .Q(n16916), .QN(n26600)
         );
  DFF_X2 avector30_reg_8__0_ ( .D(n24730), .CK(clk), .Q(n16953), .QN(n26599)
         );
  DFF_X2 avector23_reg_8__15_ ( .D(n23539), .CK(clk), .Q(n16999), .QN(n26566)
         );
  DFF_X2 avector23_reg_8__14_ ( .D(n23538), .CK(clk), .Q(n17036), .QN(n26565)
         );
  DFF_X2 avector23_reg_8__13_ ( .D(n23537), .CK(clk), .Q(n17073), .QN(n26564)
         );
  DFF_X2 avector23_reg_8__12_ ( .D(n23536), .CK(clk), .Q(n17110), .QN(n26563)
         );
  DFF_X2 avector23_reg_8__11_ ( .D(n23535), .CK(clk), .Q(n17147), .QN(n26562)
         );
  DFF_X2 avector23_reg_8__10_ ( .D(n23534), .CK(clk), .Q(n17184), .QN(n26561)
         );
  DFF_X2 avector23_reg_8__9_ ( .D(n23533), .CK(clk), .Q(n17221), .QN(n26560)
         );
  DFF_X2 avector23_reg_8__8_ ( .D(n23532), .CK(clk), .Q(n17258), .QN(n26559)
         );
  DFF_X2 avector23_reg_8__7_ ( .D(n23531), .CK(clk), .Q(n17295), .QN(n26558)
         );
  DFF_X2 avector23_reg_8__6_ ( .D(n23530), .CK(clk), .Q(n17332), .QN(n26557)
         );
  DFF_X2 avector23_reg_8__5_ ( .D(n23529), .CK(clk), .Q(n17369), .QN(n26556)
         );
  DFF_X2 avector23_reg_8__4_ ( .D(n23528), .CK(clk), .Q(n17406), .QN(n26555)
         );
  DFF_X2 avector23_reg_8__3_ ( .D(n23527), .CK(clk), .Q(n17443), .QN(n26554)
         );
  DFF_X2 avector23_reg_8__2_ ( .D(n23526), .CK(clk), .Q(n17480), .QN(n26553)
         );
  DFF_X2 avector23_reg_8__1_ ( .D(n23525), .CK(clk), .Q(n17517), .QN(n26552)
         );
  DFF_X2 avector23_reg_8__0_ ( .D(n23524), .CK(clk), .Q(n17554), .QN(n26551)
         );
  DFF_X2 avector22_reg_8__15_ ( .D(n23859), .CK(clk), .QN(n26534) );
  DFF_X2 avector22_reg_8__14_ ( .D(n23858), .CK(clk), .QN(n26533) );
  DFF_X2 avector22_reg_8__13_ ( .D(n23857), .CK(clk), .QN(n26532) );
  DFF_X2 avector22_reg_8__12_ ( .D(n23856), .CK(clk), .QN(n26531) );
  DFF_X2 avector22_reg_8__11_ ( .D(n23855), .CK(clk), .QN(n26530) );
  DFF_X2 avector22_reg_8__10_ ( .D(n23854), .CK(clk), .QN(n26529) );
  DFF_X2 avector22_reg_8__9_ ( .D(n23853), .CK(clk), .QN(n26528) );
  DFF_X2 avector22_reg_8__8_ ( .D(n23852), .CK(clk), .QN(n26527) );
  DFF_X2 avector22_reg_8__7_ ( .D(n23851), .CK(clk), .QN(n26526) );
  DFF_X2 avector22_reg_8__6_ ( .D(n23850), .CK(clk), .QN(n26525) );
  DFF_X2 avector22_reg_8__5_ ( .D(n23849), .CK(clk), .QN(n26524) );
  DFF_X2 avector22_reg_8__4_ ( .D(n23848), .CK(clk), .QN(n26523) );
  DFF_X2 avector22_reg_8__3_ ( .D(n23847), .CK(clk), .QN(n26522) );
  DFF_X2 avector22_reg_8__2_ ( .D(n23846), .CK(clk), .QN(n26521) );
  DFF_X2 avector22_reg_8__1_ ( .D(n23845), .CK(clk), .QN(n26520) );
  DFF_X2 avector22_reg_8__0_ ( .D(n23844), .CK(clk), .QN(n26519) );
  DFF_X2 avector21_reg_8__15_ ( .D(n24179), .CK(clk), .QN(n26630) );
  DFF_X2 avector21_reg_8__14_ ( .D(n24178), .CK(clk), .QN(n26629) );
  DFF_X2 avector21_reg_8__13_ ( .D(n24177), .CK(clk), .QN(n26628) );
  DFF_X2 avector21_reg_8__12_ ( .D(n24176), .CK(clk), .QN(n26627) );
  DFF_X2 avector21_reg_8__11_ ( .D(n24175), .CK(clk), .QN(n26626) );
  DFF_X2 avector21_reg_8__10_ ( .D(n24174), .CK(clk), .QN(n26625) );
  DFF_X2 avector21_reg_8__9_ ( .D(n24173), .CK(clk), .QN(n26624) );
  DFF_X2 avector21_reg_8__8_ ( .D(n24172), .CK(clk), .QN(n26623) );
  DFF_X2 avector21_reg_8__7_ ( .D(n24171), .CK(clk), .QN(n26622) );
  DFF_X2 avector21_reg_8__6_ ( .D(n24170), .CK(clk), .QN(n26621) );
  DFF_X2 avector21_reg_8__5_ ( .D(n24169), .CK(clk), .QN(n26620) );
  DFF_X2 avector21_reg_8__4_ ( .D(n24168), .CK(clk), .QN(n26619) );
  DFF_X2 avector21_reg_8__3_ ( .D(n24167), .CK(clk), .QN(n26618) );
  DFF_X2 avector21_reg_8__2_ ( .D(n24166), .CK(clk), .QN(n26617) );
  DFF_X2 avector21_reg_8__1_ ( .D(n24165), .CK(clk), .QN(n26616) );
  DFF_X2 avector21_reg_8__0_ ( .D(n24164), .CK(clk), .QN(n26615) );
  DFF_X2 avector20_reg_8__15_ ( .D(n24499), .CK(clk), .Q(n16990), .QN(n26598)
         );
  DFF_X2 avector20_reg_8__14_ ( .D(n24498), .CK(clk), .Q(n17027), .QN(n26597)
         );
  DFF_X2 avector20_reg_8__13_ ( .D(n24497), .CK(clk), .Q(n17064), .QN(n26596)
         );
  DFF_X2 avector20_reg_8__12_ ( .D(n24496), .CK(clk), .Q(n17101), .QN(n26595)
         );
  DFF_X2 avector20_reg_8__11_ ( .D(n24495), .CK(clk), .Q(n17138), .QN(n26594)
         );
  DFF_X2 avector20_reg_8__10_ ( .D(n24494), .CK(clk), .Q(n17175), .QN(n26593)
         );
  DFF_X2 avector20_reg_8__9_ ( .D(n24493), .CK(clk), .Q(n17212), .QN(n26592)
         );
  DFF_X2 avector20_reg_8__8_ ( .D(n24492), .CK(clk), .Q(n17249), .QN(n26591)
         );
  DFF_X2 avector20_reg_8__7_ ( .D(n24491), .CK(clk), .Q(n17286), .QN(n26590)
         );
  DFF_X2 avector20_reg_8__6_ ( .D(n24490), .CK(clk), .Q(n17323), .QN(n26589)
         );
  DFF_X2 avector20_reg_8__5_ ( .D(n24489), .CK(clk), .Q(n17360), .QN(n26588)
         );
  DFF_X2 avector20_reg_8__4_ ( .D(n24488), .CK(clk), .Q(n17397), .QN(n26587)
         );
  DFF_X2 avector20_reg_8__3_ ( .D(n24487), .CK(clk), .Q(n17434), .QN(n26586)
         );
  DFF_X2 avector20_reg_8__2_ ( .D(n24486), .CK(clk), .Q(n17471), .QN(n26585)
         );
  DFF_X2 avector20_reg_8__1_ ( .D(n24485), .CK(clk), .Q(n17508), .QN(n26584)
         );
  DFF_X2 avector20_reg_8__0_ ( .D(n24484), .CK(clk), .Q(n17545), .QN(n26583)
         );
  DFF_X2 avector13_reg_8__15_ ( .D(n23619), .CK(clk), .Q(n17591), .QN(n26726)
         );
  DFF_X2 avector13_reg_8__14_ ( .D(n23618), .CK(clk), .Q(n17628), .QN(n26725)
         );
  DFF_X2 avector13_reg_8__13_ ( .D(n23617), .CK(clk), .Q(n17665), .QN(n26724)
         );
  DFF_X2 avector13_reg_8__12_ ( .D(n23616), .CK(clk), .Q(n17702), .QN(n26723)
         );
  DFF_X2 avector13_reg_8__11_ ( .D(n23615), .CK(clk), .Q(n17739), .QN(n26722)
         );
  DFF_X2 avector13_reg_8__10_ ( .D(n23614), .CK(clk), .Q(n17776), .QN(n26721)
         );
  DFF_X2 avector13_reg_8__9_ ( .D(n23613), .CK(clk), .Q(n17813), .QN(n26720)
         );
  DFF_X2 avector13_reg_8__8_ ( .D(n23612), .CK(clk), .Q(n17850), .QN(n26719)
         );
  DFF_X2 avector13_reg_8__7_ ( .D(n23611), .CK(clk), .Q(n17887), .QN(n26718)
         );
  DFF_X2 avector13_reg_8__6_ ( .D(n23610), .CK(clk), .Q(n17924), .QN(n26717)
         );
  DFF_X2 avector13_reg_8__5_ ( .D(n23609), .CK(clk), .Q(n17961), .QN(n26716)
         );
  DFF_X2 avector13_reg_8__4_ ( .D(n23608), .CK(clk), .Q(n17998), .QN(n26715)
         );
  DFF_X2 avector13_reg_8__3_ ( .D(n23607), .CK(clk), .Q(n18035), .QN(n26714)
         );
  DFF_X2 avector13_reg_8__2_ ( .D(n23606), .CK(clk), .Q(n18072), .QN(n26713)
         );
  DFF_X2 avector13_reg_8__1_ ( .D(n23605), .CK(clk), .Q(n18109), .QN(n26712)
         );
  DFF_X2 avector13_reg_8__0_ ( .D(n23604), .CK(clk), .Q(n18146), .QN(n26711)
         );
  DFF_X2 avector12_reg_8__15_ ( .D(n23939), .CK(clk), .QN(n26742) );
  DFF_X2 avector12_reg_8__14_ ( .D(n23938), .CK(clk), .QN(n26741) );
  DFF_X2 avector12_reg_8__13_ ( .D(n23937), .CK(clk), .QN(n26740) );
  DFF_X2 avector12_reg_8__12_ ( .D(n23936), .CK(clk), .QN(n26739) );
  DFF_X2 avector12_reg_8__11_ ( .D(n23935), .CK(clk), .QN(n26738) );
  DFF_X2 avector12_reg_8__10_ ( .D(n23934), .CK(clk), .QN(n26737) );
  DFF_X2 avector12_reg_8__9_ ( .D(n23933), .CK(clk), .QN(n26736) );
  DFF_X2 avector12_reg_8__8_ ( .D(n23932), .CK(clk), .QN(n26735) );
  DFF_X2 avector12_reg_8__7_ ( .D(n23931), .CK(clk), .QN(n26734) );
  DFF_X2 avector12_reg_8__6_ ( .D(n23930), .CK(clk), .QN(n26733) );
  DFF_X2 avector12_reg_8__5_ ( .D(n23929), .CK(clk), .QN(n26732) );
  DFF_X2 avector12_reg_8__4_ ( .D(n23928), .CK(clk), .QN(n26731) );
  DFF_X2 avector12_reg_8__3_ ( .D(n23927), .CK(clk), .QN(n26730) );
  DFF_X2 avector12_reg_8__2_ ( .D(n23926), .CK(clk), .QN(n26729) );
  DFF_X2 avector12_reg_8__1_ ( .D(n23925), .CK(clk), .QN(n26728) );
  DFF_X2 avector12_reg_8__0_ ( .D(n23924), .CK(clk), .QN(n26727) );
  DFF_X2 avector11_reg_8__15_ ( .D(n24259), .CK(clk), .QN(n26758) );
  DFF_X2 avector11_reg_8__14_ ( .D(n24258), .CK(clk), .QN(n26757) );
  DFF_X2 avector11_reg_8__13_ ( .D(n24257), .CK(clk), .QN(n26756) );
  DFF_X2 avector11_reg_8__12_ ( .D(n24256), .CK(clk), .QN(n26755) );
  DFF_X2 avector11_reg_8__11_ ( .D(n24255), .CK(clk), .QN(n26754) );
  DFF_X2 avector11_reg_8__10_ ( .D(n24254), .CK(clk), .QN(n26753) );
  DFF_X2 avector11_reg_8__9_ ( .D(n24253), .CK(clk), .QN(n26752) );
  DFF_X2 avector11_reg_8__8_ ( .D(n24252), .CK(clk), .QN(n26751) );
  DFF_X2 avector11_reg_8__7_ ( .D(n24251), .CK(clk), .QN(n26750) );
  DFF_X2 avector11_reg_8__6_ ( .D(n24250), .CK(clk), .QN(n26749) );
  DFF_X2 avector11_reg_8__5_ ( .D(n24249), .CK(clk), .QN(n26748) );
  DFF_X2 avector11_reg_8__4_ ( .D(n24248), .CK(clk), .QN(n26747) );
  DFF_X2 avector11_reg_8__3_ ( .D(n24247), .CK(clk), .QN(n26746) );
  DFF_X2 avector11_reg_8__2_ ( .D(n24246), .CK(clk), .QN(n26745) );
  DFF_X2 avector11_reg_8__1_ ( .D(n24245), .CK(clk), .QN(n26744) );
  DFF_X2 avector11_reg_8__0_ ( .D(n24244), .CK(clk), .QN(n26743) );
  DFF_X2 avector10_reg_8__15_ ( .D(n24579), .CK(clk), .Q(n17582), .QN(n26774)
         );
  DFF_X2 avector10_reg_8__14_ ( .D(n24578), .CK(clk), .Q(n17619), .QN(n26773)
         );
  DFF_X2 avector10_reg_8__13_ ( .D(n24577), .CK(clk), .Q(n17656), .QN(n26772)
         );
  DFF_X2 avector10_reg_8__12_ ( .D(n24576), .CK(clk), .Q(n17693), .QN(n26771)
         );
  DFF_X2 avector10_reg_8__11_ ( .D(n24575), .CK(clk), .Q(n17730), .QN(n26770)
         );
  DFF_X2 avector10_reg_8__10_ ( .D(n24574), .CK(clk), .Q(n17767), .QN(n26769)
         );
  DFF_X2 avector10_reg_8__9_ ( .D(n24573), .CK(clk), .Q(n17804), .QN(n26768)
         );
  DFF_X2 avector10_reg_8__8_ ( .D(n24572), .CK(clk), .Q(n17841), .QN(n26767)
         );
  DFF_X2 avector10_reg_8__7_ ( .D(n24571), .CK(clk), .Q(n17878), .QN(n26766)
         );
  DFF_X2 avector10_reg_8__6_ ( .D(n24570), .CK(clk), .Q(n17915), .QN(n26765)
         );
  DFF_X2 avector10_reg_8__5_ ( .D(n24569), .CK(clk), .Q(n17952), .QN(n26764)
         );
  DFF_X2 avector10_reg_8__4_ ( .D(n24568), .CK(clk), .Q(n17989), .QN(n26763)
         );
  DFF_X2 avector10_reg_8__3_ ( .D(n24567), .CK(clk), .Q(n18026), .QN(n26762)
         );
  DFF_X2 avector10_reg_8__2_ ( .D(n24566), .CK(clk), .Q(n18063), .QN(n26761)
         );
  DFF_X2 avector10_reg_8__1_ ( .D(n24565), .CK(clk), .Q(n18100), .QN(n26760)
         );
  DFF_X2 avector10_reg_8__0_ ( .D(n24564), .CK(clk), .Q(n18137), .QN(n26759)
         );
  DFF_X2 avector03_reg_8__15_ ( .D(n23699), .CK(clk), .Q(n18183), .QN(n26662)
         );
  DFF_X2 avector03_reg_8__14_ ( .D(n23698), .CK(clk), .Q(n18220), .QN(n26661)
         );
  DFF_X2 avector03_reg_8__13_ ( .D(n23697), .CK(clk), .Q(n18257), .QN(n26660)
         );
  DFF_X2 avector03_reg_8__12_ ( .D(n23696), .CK(clk), .Q(n18294), .QN(n26659)
         );
  DFF_X2 avector03_reg_8__11_ ( .D(n23695), .CK(clk), .Q(n18331), .QN(n26658)
         );
  DFF_X2 avector03_reg_8__10_ ( .D(n23694), .CK(clk), .Q(n18368), .QN(n26657)
         );
  DFF_X2 avector03_reg_8__9_ ( .D(n23693), .CK(clk), .Q(n18405), .QN(n26656)
         );
  DFF_X2 avector03_reg_8__8_ ( .D(n23692), .CK(clk), .Q(n18442), .QN(n26655)
         );
  DFF_X2 avector03_reg_8__7_ ( .D(n23691), .CK(clk), .Q(n18479), .QN(n26654)
         );
  DFF_X2 avector03_reg_8__6_ ( .D(n23690), .CK(clk), .Q(n18516), .QN(n26653)
         );
  DFF_X2 avector03_reg_8__5_ ( .D(n23689), .CK(clk), .Q(n18553), .QN(n26652)
         );
  DFF_X2 avector03_reg_8__4_ ( .D(n23688), .CK(clk), .Q(n18590), .QN(n26651)
         );
  DFF_X2 avector03_reg_8__3_ ( .D(n23687), .CK(clk), .Q(n18627), .QN(n26650)
         );
  DFF_X2 avector03_reg_8__2_ ( .D(n23686), .CK(clk), .Q(n18664), .QN(n26649)
         );
  DFF_X2 avector03_reg_8__1_ ( .D(n23685), .CK(clk), .Q(n18701), .QN(n26648)
         );
  DFF_X2 avector03_reg_8__0_ ( .D(n23684), .CK(clk), .Q(n18738), .QN(n26647)
         );
  DFF_X2 avector02_reg_8__15_ ( .D(n24019), .CK(clk), .QN(n26678) );
  DFF_X2 avector02_reg_8__14_ ( .D(n24018), .CK(clk), .QN(n26677) );
  DFF_X2 avector02_reg_8__13_ ( .D(n24017), .CK(clk), .QN(n26676) );
  DFF_X2 avector02_reg_8__12_ ( .D(n24016), .CK(clk), .QN(n26675) );
  DFF_X2 avector02_reg_8__11_ ( .D(n24015), .CK(clk), .QN(n26674) );
  DFF_X2 avector02_reg_8__10_ ( .D(n24014), .CK(clk), .QN(n26673) );
  DFF_X2 avector02_reg_8__9_ ( .D(n24013), .CK(clk), .QN(n26672) );
  DFF_X2 avector02_reg_8__8_ ( .D(n24012), .CK(clk), .QN(n26671) );
  DFF_X2 avector02_reg_8__7_ ( .D(n24011), .CK(clk), .QN(n26670) );
  DFF_X2 avector02_reg_8__6_ ( .D(n24010), .CK(clk), .QN(n26669) );
  DFF_X2 avector02_reg_8__5_ ( .D(n24009), .CK(clk), .QN(n26668) );
  DFF_X2 avector02_reg_8__4_ ( .D(n24008), .CK(clk), .QN(n26667) );
  DFF_X2 avector02_reg_8__3_ ( .D(n24007), .CK(clk), .QN(n26666) );
  DFF_X2 avector02_reg_8__2_ ( .D(n24006), .CK(clk), .QN(n26665) );
  DFF_X2 avector02_reg_8__1_ ( .D(n24005), .CK(clk), .QN(n26664) );
  DFF_X2 avector02_reg_8__0_ ( .D(n24004), .CK(clk), .QN(n26663) );
  DFF_X2 avector01_reg_8__15_ ( .D(n24339), .CK(clk), .QN(n26694) );
  DFF_X2 avector01_reg_8__14_ ( .D(n24338), .CK(clk), .QN(n26693) );
  DFF_X2 avector01_reg_8__13_ ( .D(n24337), .CK(clk), .QN(n26692) );
  DFF_X2 avector01_reg_8__12_ ( .D(n24336), .CK(clk), .QN(n26691) );
  DFF_X2 avector01_reg_8__11_ ( .D(n24335), .CK(clk), .QN(n26690) );
  DFF_X2 avector01_reg_8__10_ ( .D(n24334), .CK(clk), .QN(n26689) );
  DFF_X2 avector01_reg_8__9_ ( .D(n24333), .CK(clk), .QN(n26688) );
  DFF_X2 avector01_reg_8__8_ ( .D(n24332), .CK(clk), .QN(n26687) );
  DFF_X2 avector01_reg_8__7_ ( .D(n24331), .CK(clk), .QN(n26686) );
  DFF_X2 avector01_reg_8__6_ ( .D(n24330), .CK(clk), .QN(n26685) );
  DFF_X2 avector01_reg_8__5_ ( .D(n24329), .CK(clk), .QN(n26684) );
  DFF_X2 avector01_reg_8__4_ ( .D(n24328), .CK(clk), .QN(n26683) );
  DFF_X2 avector01_reg_8__3_ ( .D(n24327), .CK(clk), .QN(n26682) );
  DFF_X2 avector01_reg_8__2_ ( .D(n24326), .CK(clk), .QN(n26681) );
  DFF_X2 avector01_reg_8__1_ ( .D(n24325), .CK(clk), .QN(n26680) );
  DFF_X2 avector01_reg_8__0_ ( .D(n24324), .CK(clk), .QN(n26679) );
  DFF_X2 avector00_reg_8__15_ ( .D(n24665), .CK(clk), .Q(n18174), .QN(n26710)
         );
  DFF_X2 avector00_reg_8__14_ ( .D(n24664), .CK(clk), .Q(n18211), .QN(n26709)
         );
  DFF_X2 avector00_reg_8__13_ ( .D(n24663), .CK(clk), .Q(n18248), .QN(n26708)
         );
  DFF_X2 avector00_reg_8__12_ ( .D(n24662), .CK(clk), .Q(n18285), .QN(n26707)
         );
  DFF_X2 avector00_reg_8__11_ ( .D(n24661), .CK(clk), .Q(n18322), .QN(n26706)
         );
  DFF_X2 avector00_reg_8__10_ ( .D(n24660), .CK(clk), .Q(n18359), .QN(n26705)
         );
  DFF_X2 avector00_reg_8__9_ ( .D(n24659), .CK(clk), .Q(n18396), .QN(n26704)
         );
  DFF_X2 avector00_reg_8__8_ ( .D(n24658), .CK(clk), .Q(n18433), .QN(n26703)
         );
  DFF_X2 avector00_reg_8__7_ ( .D(n24657), .CK(clk), .Q(n18470), .QN(n26702)
         );
  DFF_X2 avector00_reg_8__6_ ( .D(n24656), .CK(clk), .Q(n18507), .QN(n26701)
         );
  DFF_X2 avector00_reg_8__5_ ( .D(n24655), .CK(clk), .Q(n18544), .QN(n26700)
         );
  DFF_X2 avector00_reg_8__4_ ( .D(n24654), .CK(clk), .Q(n18581), .QN(n26699)
         );
  DFF_X2 avector00_reg_8__3_ ( .D(n24653), .CK(clk), .Q(n18618), .QN(n26698)
         );
  DFF_X2 avector00_reg_8__2_ ( .D(n24652), .CK(clk), .Q(n18655), .QN(n26697)
         );
  DFF_X2 avector00_reg_8__1_ ( .D(n24651), .CK(clk), .Q(n18692), .QN(n26696)
         );
  DFF_X2 avector00_reg_8__0_ ( .D(n24650), .CK(clk), .Q(n18729), .QN(n26695)
         );
  DFF_X2 avector33_reg_7__15_ ( .D(n23795), .CK(clk), .QN(n27606) );
  DFF_X2 avector33_reg_7__14_ ( .D(n23794), .CK(clk), .QN(n27605) );
  DFF_X2 avector33_reg_7__13_ ( .D(n23793), .CK(clk), .QN(n27604) );
  DFF_X2 avector33_reg_7__12_ ( .D(n23792), .CK(clk), .QN(n27603) );
  DFF_X2 avector33_reg_7__11_ ( .D(n23791), .CK(clk), .QN(n27602) );
  DFF_X2 avector33_reg_7__10_ ( .D(n23790), .CK(clk), .QN(n27601) );
  DFF_X2 avector33_reg_7__9_ ( .D(n23789), .CK(clk), .QN(n27600) );
  DFF_X2 avector33_reg_7__8_ ( .D(n23788), .CK(clk), .QN(n27599) );
  DFF_X2 avector33_reg_7__7_ ( .D(n23787), .CK(clk), .QN(n27598) );
  DFF_X2 avector33_reg_7__6_ ( .D(n23786), .CK(clk), .QN(n27597) );
  DFF_X2 avector33_reg_7__5_ ( .D(n23785), .CK(clk), .QN(n27596) );
  DFF_X2 avector33_reg_7__4_ ( .D(n23784), .CK(clk), .QN(n27595) );
  DFF_X2 avector33_reg_7__3_ ( .D(n23783), .CK(clk), .QN(n27594) );
  DFF_X2 avector33_reg_7__2_ ( .D(n23782), .CK(clk), .QN(n27593) );
  DFF_X2 avector33_reg_7__1_ ( .D(n23781), .CK(clk), .QN(n27592) );
  DFF_X2 avector33_reg_7__0_ ( .D(n23780), .CK(clk), .QN(n27591) );
  DFF_X2 avector33_reg_6__15_ ( .D(n23811), .CK(clk), .QN(n26838) );
  DFF_X2 avector33_reg_6__14_ ( .D(n23810), .CK(clk), .QN(n26837) );
  DFF_X2 avector33_reg_6__13_ ( .D(n23809), .CK(clk), .QN(n26836) );
  DFF_X2 avector33_reg_6__12_ ( .D(n23808), .CK(clk), .QN(n26835) );
  DFF_X2 avector33_reg_6__11_ ( .D(n23807), .CK(clk), .QN(n26834) );
  DFF_X2 avector33_reg_6__10_ ( .D(n23806), .CK(clk), .QN(n26833) );
  DFF_X2 avector33_reg_6__9_ ( .D(n23805), .CK(clk), .QN(n26832) );
  DFF_X2 avector33_reg_6__8_ ( .D(n23804), .CK(clk), .QN(n26831) );
  DFF_X2 avector33_reg_6__7_ ( .D(n23803), .CK(clk), .QN(n26830) );
  DFF_X2 avector33_reg_6__6_ ( .D(n23802), .CK(clk), .QN(n26829) );
  DFF_X2 avector33_reg_6__5_ ( .D(n23801), .CK(clk), .QN(n26828) );
  DFF_X2 avector33_reg_6__4_ ( .D(n23800), .CK(clk), .QN(n26827) );
  DFF_X2 avector33_reg_6__3_ ( .D(n23799), .CK(clk), .QN(n26826) );
  DFF_X2 avector33_reg_6__2_ ( .D(n23798), .CK(clk), .QN(n26825) );
  DFF_X2 avector33_reg_6__1_ ( .D(n23797), .CK(clk), .QN(n26824) );
  DFF_X2 avector33_reg_6__0_ ( .D(n23796), .CK(clk), .QN(n26823) );
  DFF_X2 avector33_reg_1__15_ ( .D(n23827), .CK(clk), .Q(n16402), .QN(n27094)
         );
  DFF_X2 avector33_reg_1__14_ ( .D(n23826), .CK(clk), .Q(n16439), .QN(n27093)
         );
  DFF_X2 avector33_reg_1__13_ ( .D(n23825), .CK(clk), .Q(n16476), .QN(n27092)
         );
  DFF_X2 avector33_reg_1__12_ ( .D(n23824), .CK(clk), .Q(n16513), .QN(n27091)
         );
  DFF_X2 avector33_reg_1__11_ ( .D(n23823), .CK(clk), .Q(n16550), .QN(n27090)
         );
  DFF_X2 avector33_reg_1__10_ ( .D(n23822), .CK(clk), .Q(n16587), .QN(n27089)
         );
  DFF_X2 avector33_reg_1__9_ ( .D(n23821), .CK(clk), .Q(n16624), .QN(n27088)
         );
  DFF_X2 avector33_reg_1__8_ ( .D(n23820), .CK(clk), .Q(n16661), .QN(n27087)
         );
  DFF_X2 avector33_reg_1__7_ ( .D(n23819), .CK(clk), .Q(n16698), .QN(n27086)
         );
  DFF_X2 avector33_reg_1__6_ ( .D(n23818), .CK(clk), .Q(n16735), .QN(n27085)
         );
  DFF_X2 avector33_reg_1__5_ ( .D(n23817), .CK(clk), .Q(n16772), .QN(n27084)
         );
  DFF_X2 avector33_reg_1__4_ ( .D(n23816), .CK(clk), .Q(n16809), .QN(n27083)
         );
  DFF_X2 avector33_reg_1__3_ ( .D(n23815), .CK(clk), .Q(n16846), .QN(n27082)
         );
  DFF_X2 avector33_reg_1__2_ ( .D(n23814), .CK(clk), .Q(n16883), .QN(n27081)
         );
  DFF_X2 avector33_reg_1__1_ ( .D(n23813), .CK(clk), .Q(n16920), .QN(n27080)
         );
  DFF_X2 avector33_reg_1__0_ ( .D(n23812), .CK(clk), .Q(n16957), .QN(n27079)
         );
  DFF_X2 avector33_reg_0__15_ ( .D(n23843), .CK(clk), .Q(n16403), .QN(n27350)
         );
  DFF_X2 avector33_reg_0__14_ ( .D(n23842), .CK(clk), .Q(n16440), .QN(n27349)
         );
  DFF_X2 avector33_reg_0__13_ ( .D(n23841), .CK(clk), .Q(n16477), .QN(n27348)
         );
  DFF_X2 avector33_reg_0__12_ ( .D(n23840), .CK(clk), .Q(n16514), .QN(n27347)
         );
  DFF_X2 avector33_reg_0__11_ ( .D(n23839), .CK(clk), .Q(n16551), .QN(n27346)
         );
  DFF_X2 avector33_reg_0__10_ ( .D(n23838), .CK(clk), .Q(n16588), .QN(n27345)
         );
  DFF_X2 avector33_reg_0__9_ ( .D(n23837), .CK(clk), .Q(n16625), .QN(n27344)
         );
  DFF_X2 avector33_reg_0__8_ ( .D(n23836), .CK(clk), .Q(n16662), .QN(n27343)
         );
  DFF_X2 avector33_reg_0__7_ ( .D(n23835), .CK(clk), .Q(n16699), .QN(n27342)
         );
  DFF_X2 avector33_reg_0__6_ ( .D(n23834), .CK(clk), .Q(n16736), .QN(n27341)
         );
  DFF_X2 avector33_reg_0__5_ ( .D(n23833), .CK(clk), .Q(n16773), .QN(n27340)
         );
  DFF_X2 avector33_reg_0__4_ ( .D(n23832), .CK(clk), .Q(n16810), .QN(n27339)
         );
  DFF_X2 avector33_reg_0__3_ ( .D(n23831), .CK(clk), .Q(n16847), .QN(n27338)
         );
  DFF_X2 avector33_reg_0__2_ ( .D(n23830), .CK(clk), .Q(n16884), .QN(n27337)
         );
  DFF_X2 avector33_reg_0__1_ ( .D(n23829), .CK(clk), .Q(n16921), .QN(n27336)
         );
  DFF_X2 avector33_reg_0__0_ ( .D(n23828), .CK(clk), .Q(n16958), .QN(n27335)
         );
  DFF_X2 avector32_reg_7__15_ ( .D(n24115), .CK(clk), .Q(n16381), .QN(n27670)
         );
  DFF_X2 avector32_reg_7__14_ ( .D(n24114), .CK(clk), .Q(n16418), .QN(n27669)
         );
  DFF_X2 avector32_reg_7__13_ ( .D(n24113), .CK(clk), .Q(n16455), .QN(n27668)
         );
  DFF_X2 avector32_reg_7__12_ ( .D(n24112), .CK(clk), .Q(n16492), .QN(n27667)
         );
  DFF_X2 avector32_reg_7__11_ ( .D(n24111), .CK(clk), .Q(n16529), .QN(n27666)
         );
  DFF_X2 avector32_reg_7__10_ ( .D(n24110), .CK(clk), .Q(n16566), .QN(n27665)
         );
  DFF_X2 avector32_reg_7__9_ ( .D(n24109), .CK(clk), .Q(n16603), .QN(n27664)
         );
  DFF_X2 avector32_reg_7__8_ ( .D(n24108), .CK(clk), .Q(n16640), .QN(n27663)
         );
  DFF_X2 avector32_reg_7__7_ ( .D(n24107), .CK(clk), .Q(n16677), .QN(n27662)
         );
  DFF_X2 avector32_reg_7__6_ ( .D(n24106), .CK(clk), .Q(n16714), .QN(n27661)
         );
  DFF_X2 avector32_reg_7__5_ ( .D(n24105), .CK(clk), .Q(n16751), .QN(n27660)
         );
  DFF_X2 avector32_reg_7__4_ ( .D(n24104), .CK(clk), .Q(n16788), .QN(n27659)
         );
  DFF_X2 avector32_reg_7__3_ ( .D(n24103), .CK(clk), .Q(n16825), .QN(n27658)
         );
  DFF_X2 avector32_reg_7__2_ ( .D(n24102), .CK(clk), .Q(n16862), .QN(n27657)
         );
  DFF_X2 avector32_reg_7__1_ ( .D(n24101), .CK(clk), .Q(n16899), .QN(n27656)
         );
  DFF_X2 avector32_reg_7__0_ ( .D(n24100), .CK(clk), .Q(n16936), .QN(n27655)
         );
  DFF_X2 avector32_reg_6__15_ ( .D(n24131), .CK(clk), .Q(n16379), .QN(n26902)
         );
  DFF_X2 avector32_reg_6__14_ ( .D(n24130), .CK(clk), .Q(n16416), .QN(n26901)
         );
  DFF_X2 avector32_reg_6__13_ ( .D(n24129), .CK(clk), .Q(n16453), .QN(n26900)
         );
  DFF_X2 avector32_reg_6__12_ ( .D(n24128), .CK(clk), .Q(n16490), .QN(n26899)
         );
  DFF_X2 avector32_reg_6__11_ ( .D(n24127), .CK(clk), .Q(n16527), .QN(n26898)
         );
  DFF_X2 avector32_reg_6__10_ ( .D(n24126), .CK(clk), .Q(n16564), .QN(n26897)
         );
  DFF_X2 avector32_reg_6__9_ ( .D(n24125), .CK(clk), .Q(n16601), .QN(n26896)
         );
  DFF_X2 avector32_reg_6__8_ ( .D(n24124), .CK(clk), .Q(n16638), .QN(n26895)
         );
  DFF_X2 avector32_reg_6__7_ ( .D(n24123), .CK(clk), .Q(n16675), .QN(n26894)
         );
  DFF_X2 avector32_reg_6__6_ ( .D(n24122), .CK(clk), .Q(n16712), .QN(n26893)
         );
  DFF_X2 avector32_reg_6__5_ ( .D(n24121), .CK(clk), .Q(n16749), .QN(n26892)
         );
  DFF_X2 avector32_reg_6__4_ ( .D(n24120), .CK(clk), .Q(n16786), .QN(n26891)
         );
  DFF_X2 avector32_reg_6__3_ ( .D(n24119), .CK(clk), .Q(n16823), .QN(n26890)
         );
  DFF_X2 avector32_reg_6__2_ ( .D(n24118), .CK(clk), .Q(n16860), .QN(n26889)
         );
  DFF_X2 avector32_reg_6__1_ ( .D(n24117), .CK(clk), .Q(n16897), .QN(n26888)
         );
  DFF_X2 avector32_reg_6__0_ ( .D(n24116), .CK(clk), .Q(n16934), .QN(n26887)
         );
  DFF_X2 avector32_reg_1__15_ ( .D(n24147), .CK(clk), .QN(n27158) );
  DFF_X2 avector32_reg_1__14_ ( .D(n24146), .CK(clk), .QN(n27157) );
  DFF_X2 avector32_reg_1__13_ ( .D(n24145), .CK(clk), .QN(n27156) );
  DFF_X2 avector32_reg_1__12_ ( .D(n24144), .CK(clk), .QN(n27155) );
  DFF_X2 avector32_reg_1__11_ ( .D(n24143), .CK(clk), .QN(n27154) );
  DFF_X2 avector32_reg_1__10_ ( .D(n24142), .CK(clk), .QN(n27153) );
  DFF_X2 avector32_reg_1__9_ ( .D(n24141), .CK(clk), .QN(n27152) );
  DFF_X2 avector32_reg_1__8_ ( .D(n24140), .CK(clk), .QN(n27151) );
  DFF_X2 avector32_reg_1__7_ ( .D(n24139), .CK(clk), .QN(n27150) );
  DFF_X2 avector32_reg_1__6_ ( .D(n24138), .CK(clk), .QN(n27149) );
  DFF_X2 avector32_reg_1__5_ ( .D(n24137), .CK(clk), .QN(n27148) );
  DFF_X2 avector32_reg_1__4_ ( .D(n24136), .CK(clk), .QN(n27147) );
  DFF_X2 avector32_reg_1__3_ ( .D(n24135), .CK(clk), .QN(n27146) );
  DFF_X2 avector32_reg_1__2_ ( .D(n24134), .CK(clk), .QN(n27145) );
  DFF_X2 avector32_reg_1__1_ ( .D(n24133), .CK(clk), .QN(n27144) );
  DFF_X2 avector32_reg_1__0_ ( .D(n24132), .CK(clk), .QN(n27143) );
  DFF_X2 avector32_reg_0__15_ ( .D(n24163), .CK(clk), .QN(n27414) );
  DFF_X2 avector32_reg_0__14_ ( .D(n24162), .CK(clk), .QN(n27413) );
  DFF_X2 avector32_reg_0__13_ ( .D(n24161), .CK(clk), .QN(n27412) );
  DFF_X2 avector32_reg_0__12_ ( .D(n24160), .CK(clk), .QN(n27411) );
  DFF_X2 avector32_reg_0__11_ ( .D(n24159), .CK(clk), .QN(n27410) );
  DFF_X2 avector32_reg_0__10_ ( .D(n24158), .CK(clk), .QN(n27409) );
  DFF_X2 avector32_reg_0__9_ ( .D(n24157), .CK(clk), .QN(n27408) );
  DFF_X2 avector32_reg_0__8_ ( .D(n24156), .CK(clk), .QN(n27407) );
  DFF_X2 avector32_reg_0__7_ ( .D(n24155), .CK(clk), .QN(n27406) );
  DFF_X2 avector32_reg_0__6_ ( .D(n24154), .CK(clk), .QN(n27405) );
  DFF_X2 avector32_reg_0__5_ ( .D(n24153), .CK(clk), .QN(n27404) );
  DFF_X2 avector32_reg_0__4_ ( .D(n24152), .CK(clk), .QN(n27403) );
  DFF_X2 avector32_reg_0__3_ ( .D(n24151), .CK(clk), .QN(n27402) );
  DFF_X2 avector32_reg_0__2_ ( .D(n24150), .CK(clk), .QN(n27401) );
  DFF_X2 avector32_reg_0__1_ ( .D(n24149), .CK(clk), .QN(n27400) );
  DFF_X2 avector32_reg_0__0_ ( .D(n24148), .CK(clk), .QN(n27399) );
  DFF_X2 avector31_reg_7__15_ ( .D(n24435), .CK(clk), .Q(n16390), .QN(n27734)
         );
  DFF_X2 avector31_reg_7__14_ ( .D(n24434), .CK(clk), .Q(n16427), .QN(n27733)
         );
  DFF_X2 avector31_reg_7__13_ ( .D(n24433), .CK(clk), .Q(n16464), .QN(n27732)
         );
  DFF_X2 avector31_reg_7__12_ ( .D(n24432), .CK(clk), .Q(n16501), .QN(n27731)
         );
  DFF_X2 avector31_reg_7__11_ ( .D(n24431), .CK(clk), .Q(n16538), .QN(n27730)
         );
  DFF_X2 avector31_reg_7__10_ ( .D(n24430), .CK(clk), .Q(n16575), .QN(n27729)
         );
  DFF_X2 avector31_reg_7__9_ ( .D(n24429), .CK(clk), .Q(n16612), .QN(n27728)
         );
  DFF_X2 avector31_reg_7__8_ ( .D(n24428), .CK(clk), .Q(n16649), .QN(n27727)
         );
  DFF_X2 avector31_reg_7__7_ ( .D(n24427), .CK(clk), .Q(n16686), .QN(n27726)
         );
  DFF_X2 avector31_reg_7__6_ ( .D(n24426), .CK(clk), .Q(n16723), .QN(n27725)
         );
  DFF_X2 avector31_reg_7__5_ ( .D(n24425), .CK(clk), .Q(n16760), .QN(n27724)
         );
  DFF_X2 avector31_reg_7__4_ ( .D(n24424), .CK(clk), .Q(n16797), .QN(n27723)
         );
  DFF_X2 avector31_reg_7__3_ ( .D(n24423), .CK(clk), .Q(n16834), .QN(n27722)
         );
  DFF_X2 avector31_reg_7__2_ ( .D(n24422), .CK(clk), .Q(n16871), .QN(n27721)
         );
  DFF_X2 avector31_reg_7__1_ ( .D(n24421), .CK(clk), .Q(n16908), .QN(n27720)
         );
  DFF_X2 avector31_reg_7__0_ ( .D(n24420), .CK(clk), .Q(n16945), .QN(n27719)
         );
  DFF_X2 avector31_reg_6__15_ ( .D(n24451), .CK(clk), .QN(n26966) );
  DFF_X2 avector31_reg_6__14_ ( .D(n24450), .CK(clk), .QN(n26965) );
  DFF_X2 avector31_reg_6__13_ ( .D(n24449), .CK(clk), .QN(n26964) );
  DFF_X2 avector31_reg_6__12_ ( .D(n24448), .CK(clk), .QN(n26963) );
  DFF_X2 avector31_reg_6__11_ ( .D(n24447), .CK(clk), .QN(n26962) );
  DFF_X2 avector31_reg_6__10_ ( .D(n24446), .CK(clk), .QN(n26961) );
  DFF_X2 avector31_reg_6__9_ ( .D(n24445), .CK(clk), .QN(n26960) );
  DFF_X2 avector31_reg_6__8_ ( .D(n24444), .CK(clk), .QN(n26959) );
  DFF_X2 avector31_reg_6__7_ ( .D(n24443), .CK(clk), .QN(n26958) );
  DFF_X2 avector31_reg_6__6_ ( .D(n24442), .CK(clk), .QN(n26957) );
  DFF_X2 avector31_reg_6__5_ ( .D(n24441), .CK(clk), .QN(n26956) );
  DFF_X2 avector31_reg_6__4_ ( .D(n24440), .CK(clk), .QN(n26955) );
  DFF_X2 avector31_reg_6__3_ ( .D(n24439), .CK(clk), .QN(n26954) );
  DFF_X2 avector31_reg_6__2_ ( .D(n24438), .CK(clk), .QN(n26953) );
  DFF_X2 avector31_reg_6__1_ ( .D(n24437), .CK(clk), .QN(n26952) );
  DFF_X2 avector31_reg_6__0_ ( .D(n24436), .CK(clk), .QN(n26951) );
  DFF_X2 avector31_reg_1__15_ ( .D(n24467), .CK(clk), .QN(n27222) );
  DFF_X2 avector31_reg_1__14_ ( .D(n24466), .CK(clk), .QN(n27221) );
  DFF_X2 avector31_reg_1__13_ ( .D(n24465), .CK(clk), .QN(n27220) );
  DFF_X2 avector31_reg_1__12_ ( .D(n24464), .CK(clk), .QN(n27219) );
  DFF_X2 avector31_reg_1__11_ ( .D(n24463), .CK(clk), .QN(n27218) );
  DFF_X2 avector31_reg_1__10_ ( .D(n24462), .CK(clk), .QN(n27217) );
  DFF_X2 avector31_reg_1__9_ ( .D(n24461), .CK(clk), .QN(n27216) );
  DFF_X2 avector31_reg_1__8_ ( .D(n24460), .CK(clk), .QN(n27215) );
  DFF_X2 avector31_reg_1__7_ ( .D(n24459), .CK(clk), .QN(n27214) );
  DFF_X2 avector31_reg_1__6_ ( .D(n24458), .CK(clk), .QN(n27213) );
  DFF_X2 avector31_reg_1__5_ ( .D(n24457), .CK(clk), .QN(n27212) );
  DFF_X2 avector31_reg_1__4_ ( .D(n24456), .CK(clk), .QN(n27211) );
  DFF_X2 avector31_reg_1__3_ ( .D(n24455), .CK(clk), .QN(n27210) );
  DFF_X2 avector31_reg_1__2_ ( .D(n24454), .CK(clk), .QN(n27209) );
  DFF_X2 avector31_reg_1__1_ ( .D(n24453), .CK(clk), .QN(n27208) );
  DFF_X2 avector31_reg_1__0_ ( .D(n24452), .CK(clk), .QN(n27207) );
  DFF_X2 avector31_reg_0__15_ ( .D(n24483), .CK(clk), .QN(n27478) );
  DFF_X2 avector31_reg_0__14_ ( .D(n24482), .CK(clk), .QN(n27477) );
  DFF_X2 avector31_reg_0__13_ ( .D(n24481), .CK(clk), .QN(n27476) );
  DFF_X2 avector31_reg_0__12_ ( .D(n24480), .CK(clk), .QN(n27475) );
  DFF_X2 avector31_reg_0__11_ ( .D(n24479), .CK(clk), .QN(n27474) );
  DFF_X2 avector31_reg_0__10_ ( .D(n24478), .CK(clk), .QN(n27473) );
  DFF_X2 avector31_reg_0__9_ ( .D(n24477), .CK(clk), .QN(n27472) );
  DFF_X2 avector31_reg_0__8_ ( .D(n24476), .CK(clk), .QN(n27471) );
  DFF_X2 avector31_reg_0__7_ ( .D(n24475), .CK(clk), .QN(n27470) );
  DFF_X2 avector31_reg_0__6_ ( .D(n24474), .CK(clk), .QN(n27469) );
  DFF_X2 avector31_reg_0__5_ ( .D(n24473), .CK(clk), .QN(n27468) );
  DFF_X2 avector31_reg_0__4_ ( .D(n24472), .CK(clk), .QN(n27467) );
  DFF_X2 avector31_reg_0__3_ ( .D(n24471), .CK(clk), .QN(n27466) );
  DFF_X2 avector31_reg_0__2_ ( .D(n24470), .CK(clk), .QN(n27465) );
  DFF_X2 avector31_reg_0__1_ ( .D(n24469), .CK(clk), .QN(n27464) );
  DFF_X2 avector31_reg_0__0_ ( .D(n24468), .CK(clk), .QN(n27463) );
  DFF_X2 avector30_reg_7__15_ ( .D(n24761), .CK(clk), .QN(n27798) );
  DFF_X2 avector30_reg_7__14_ ( .D(n24760), .CK(clk), .QN(n27797) );
  DFF_X2 avector30_reg_7__13_ ( .D(n24759), .CK(clk), .QN(n27796) );
  DFF_X2 avector30_reg_7__12_ ( .D(n24758), .CK(clk), .QN(n27795) );
  DFF_X2 avector30_reg_7__11_ ( .D(n24757), .CK(clk), .QN(n27794) );
  DFF_X2 avector30_reg_7__10_ ( .D(n24756), .CK(clk), .QN(n27793) );
  DFF_X2 avector30_reg_7__9_ ( .D(n24755), .CK(clk), .QN(n27792) );
  DFF_X2 avector30_reg_7__8_ ( .D(n24754), .CK(clk), .QN(n27791) );
  DFF_X2 avector30_reg_7__7_ ( .D(n24753), .CK(clk), .QN(n27790) );
  DFF_X2 avector30_reg_7__6_ ( .D(n24752), .CK(clk), .QN(n27789) );
  DFF_X2 avector30_reg_7__5_ ( .D(n24751), .CK(clk), .QN(n27788) );
  DFF_X2 avector30_reg_7__4_ ( .D(n24750), .CK(clk), .QN(n27787) );
  DFF_X2 avector30_reg_7__3_ ( .D(n24749), .CK(clk), .QN(n27786) );
  DFF_X2 avector30_reg_7__2_ ( .D(n24748), .CK(clk), .QN(n27785) );
  DFF_X2 avector30_reg_7__1_ ( .D(n24747), .CK(clk), .QN(n27784) );
  DFF_X2 avector30_reg_7__0_ ( .D(n24746), .CK(clk), .QN(n27783) );
  DFF_X2 avector30_reg_6__15_ ( .D(n24777), .CK(clk), .QN(n27030) );
  DFF_X2 avector30_reg_6__14_ ( .D(n24776), .CK(clk), .QN(n27029) );
  DFF_X2 avector30_reg_6__13_ ( .D(n24775), .CK(clk), .QN(n27028) );
  DFF_X2 avector30_reg_6__12_ ( .D(n24774), .CK(clk), .QN(n27027) );
  DFF_X2 avector30_reg_6__11_ ( .D(n24773), .CK(clk), .QN(n27026) );
  DFF_X2 avector30_reg_6__10_ ( .D(n24772), .CK(clk), .QN(n27025) );
  DFF_X2 avector30_reg_6__9_ ( .D(n24771), .CK(clk), .QN(n27024) );
  DFF_X2 avector30_reg_6__8_ ( .D(n24770), .CK(clk), .QN(n27023) );
  DFF_X2 avector30_reg_6__7_ ( .D(n24769), .CK(clk), .QN(n27022) );
  DFF_X2 avector30_reg_6__6_ ( .D(n24768), .CK(clk), .QN(n27021) );
  DFF_X2 avector30_reg_6__5_ ( .D(n24767), .CK(clk), .QN(n27020) );
  DFF_X2 avector30_reg_6__4_ ( .D(n24766), .CK(clk), .QN(n27019) );
  DFF_X2 avector30_reg_6__3_ ( .D(n24765), .CK(clk), .QN(n27018) );
  DFF_X2 avector30_reg_6__2_ ( .D(n24764), .CK(clk), .QN(n27017) );
  DFF_X2 avector30_reg_6__1_ ( .D(n24763), .CK(clk), .QN(n27016) );
  DFF_X2 avector30_reg_6__0_ ( .D(n24762), .CK(clk), .QN(n27015) );
  DFF_X2 avector30_reg_1__15_ ( .D(n24793), .CK(clk), .Q(n16393), .QN(n27286)
         );
  DFF_X2 avector30_reg_1__14_ ( .D(n24792), .CK(clk), .Q(n16430), .QN(n27285)
         );
  DFF_X2 avector30_reg_1__13_ ( .D(n24791), .CK(clk), .Q(n16467), .QN(n27284)
         );
  DFF_X2 avector30_reg_1__12_ ( .D(n24790), .CK(clk), .Q(n16504), .QN(n27283)
         );
  DFF_X2 avector30_reg_1__11_ ( .D(n24789), .CK(clk), .Q(n16541), .QN(n27282)
         );
  DFF_X2 avector30_reg_1__10_ ( .D(n24788), .CK(clk), .Q(n16578), .QN(n27281)
         );
  DFF_X2 avector30_reg_1__9_ ( .D(n24787), .CK(clk), .Q(n16615), .QN(n27280)
         );
  DFF_X2 avector30_reg_1__8_ ( .D(n24786), .CK(clk), .Q(n16652), .QN(n27279)
         );
  DFF_X2 avector30_reg_1__7_ ( .D(n24785), .CK(clk), .Q(n16689), .QN(n27278)
         );
  DFF_X2 avector30_reg_1__6_ ( .D(n24784), .CK(clk), .Q(n16726), .QN(n27277)
         );
  DFF_X2 avector30_reg_1__5_ ( .D(n24783), .CK(clk), .Q(n16763), .QN(n27276)
         );
  DFF_X2 avector30_reg_1__4_ ( .D(n24782), .CK(clk), .Q(n16800), .QN(n27275)
         );
  DFF_X2 avector30_reg_1__3_ ( .D(n24781), .CK(clk), .Q(n16837), .QN(n27274)
         );
  DFF_X2 avector30_reg_1__2_ ( .D(n24780), .CK(clk), .Q(n16874), .QN(n27273)
         );
  DFF_X2 avector30_reg_1__1_ ( .D(n24779), .CK(clk), .Q(n16911), .QN(n27272)
         );
  DFF_X2 avector30_reg_1__0_ ( .D(n24778), .CK(clk), .Q(n16948), .QN(n27271)
         );
  DFF_X2 avector23_reg_7__15_ ( .D(n23555), .CK(clk), .QN(n27558) );
  DFF_X2 avector23_reg_7__14_ ( .D(n23554), .CK(clk), .QN(n27557) );
  DFF_X2 avector23_reg_7__13_ ( .D(n23553), .CK(clk), .QN(n27556) );
  DFF_X2 avector23_reg_7__12_ ( .D(n23552), .CK(clk), .QN(n27555) );
  DFF_X2 avector23_reg_7__11_ ( .D(n23551), .CK(clk), .QN(n27554) );
  DFF_X2 avector23_reg_7__10_ ( .D(n23550), .CK(clk), .QN(n27553) );
  DFF_X2 avector23_reg_7__9_ ( .D(n23549), .CK(clk), .QN(n27552) );
  DFF_X2 avector23_reg_7__8_ ( .D(n23548), .CK(clk), .QN(n27551) );
  DFF_X2 avector23_reg_7__7_ ( .D(n23547), .CK(clk), .QN(n27550) );
  DFF_X2 avector23_reg_7__6_ ( .D(n23546), .CK(clk), .QN(n27549) );
  DFF_X2 avector23_reg_7__5_ ( .D(n23545), .CK(clk), .QN(n27548) );
  DFF_X2 avector23_reg_7__4_ ( .D(n23544), .CK(clk), .QN(n27547) );
  DFF_X2 avector23_reg_7__3_ ( .D(n23543), .CK(clk), .QN(n27546) );
  DFF_X2 avector23_reg_7__2_ ( .D(n23542), .CK(clk), .QN(n27545) );
  DFF_X2 avector23_reg_7__1_ ( .D(n23541), .CK(clk), .QN(n27544) );
  DFF_X2 avector23_reg_7__0_ ( .D(n23540), .CK(clk), .QN(n27543) );
  DFF_X2 avector23_reg_6__15_ ( .D(n23571), .CK(clk), .QN(n26790) );
  DFF_X2 avector23_reg_6__14_ ( .D(n23570), .CK(clk), .QN(n26789) );
  DFF_X2 avector23_reg_6__13_ ( .D(n23569), .CK(clk), .QN(n26788) );
  DFF_X2 avector23_reg_6__12_ ( .D(n23568), .CK(clk), .QN(n26787) );
  DFF_X2 avector23_reg_6__11_ ( .D(n23567), .CK(clk), .QN(n26786) );
  DFF_X2 avector23_reg_6__10_ ( .D(n23566), .CK(clk), .QN(n26785) );
  DFF_X2 avector23_reg_6__9_ ( .D(n23565), .CK(clk), .QN(n26784) );
  DFF_X2 avector23_reg_6__8_ ( .D(n23564), .CK(clk), .QN(n26783) );
  DFF_X2 avector23_reg_6__7_ ( .D(n23563), .CK(clk), .QN(n26782) );
  DFF_X2 avector23_reg_6__6_ ( .D(n23562), .CK(clk), .QN(n26781) );
  DFF_X2 avector23_reg_6__5_ ( .D(n23561), .CK(clk), .QN(n26780) );
  DFF_X2 avector23_reg_6__4_ ( .D(n23560), .CK(clk), .QN(n26779) );
  DFF_X2 avector23_reg_6__3_ ( .D(n23559), .CK(clk), .QN(n26778) );
  DFF_X2 avector23_reg_6__2_ ( .D(n23558), .CK(clk), .QN(n26777) );
  DFF_X2 avector23_reg_6__1_ ( .D(n23557), .CK(clk), .QN(n26776) );
  DFF_X2 avector23_reg_6__0_ ( .D(n23556), .CK(clk), .QN(n26775) );
  DFF_X2 avector23_reg_1__15_ ( .D(n23587), .CK(clk), .Q(n16994), .QN(n27046)
         );
  DFF_X2 avector23_reg_1__14_ ( .D(n23586), .CK(clk), .Q(n17031), .QN(n27045)
         );
  DFF_X2 avector23_reg_1__13_ ( .D(n23585), .CK(clk), .Q(n17068), .QN(n27044)
         );
  DFF_X2 avector23_reg_1__12_ ( .D(n23584), .CK(clk), .Q(n17105), .QN(n27043)
         );
  DFF_X2 avector23_reg_1__11_ ( .D(n23583), .CK(clk), .Q(n17142), .QN(n27042)
         );
  DFF_X2 avector23_reg_1__10_ ( .D(n23582), .CK(clk), .Q(n17179), .QN(n27041)
         );
  DFF_X2 avector23_reg_1__9_ ( .D(n23581), .CK(clk), .Q(n17216), .QN(n27040)
         );
  DFF_X2 avector23_reg_1__8_ ( .D(n23580), .CK(clk), .Q(n17253), .QN(n27039)
         );
  DFF_X2 avector23_reg_1__7_ ( .D(n23579), .CK(clk), .Q(n17290), .QN(n27038)
         );
  DFF_X2 avector23_reg_1__6_ ( .D(n23578), .CK(clk), .Q(n17327), .QN(n27037)
         );
  DFF_X2 avector23_reg_1__5_ ( .D(n23577), .CK(clk), .Q(n17364), .QN(n27036)
         );
  DFF_X2 avector23_reg_1__4_ ( .D(n23576), .CK(clk), .Q(n17401), .QN(n27035)
         );
  DFF_X2 avector23_reg_1__3_ ( .D(n23575), .CK(clk), .Q(n17438), .QN(n27034)
         );
  DFF_X2 avector23_reg_1__2_ ( .D(n23574), .CK(clk), .Q(n17475), .QN(n27033)
         );
  DFF_X2 avector23_reg_1__1_ ( .D(n23573), .CK(clk), .Q(n17512), .QN(n27032)
         );
  DFF_X2 avector23_reg_1__0_ ( .D(n23572), .CK(clk), .Q(n17549), .QN(n27031)
         );
  DFF_X2 avector23_reg_0__15_ ( .D(n23603), .CK(clk), .Q(n16995), .QN(n27302)
         );
  DFF_X2 avector23_reg_0__14_ ( .D(n23602), .CK(clk), .Q(n17032), .QN(n27301)
         );
  DFF_X2 avector23_reg_0__13_ ( .D(n23601), .CK(clk), .Q(n17069), .QN(n27300)
         );
  DFF_X2 avector23_reg_0__12_ ( .D(n23600), .CK(clk), .Q(n17106), .QN(n27299)
         );
  DFF_X2 avector23_reg_0__11_ ( .D(n23599), .CK(clk), .Q(n17143), .QN(n27298)
         );
  DFF_X2 avector23_reg_0__10_ ( .D(n23598), .CK(clk), .Q(n17180), .QN(n27297)
         );
  DFF_X2 avector23_reg_0__9_ ( .D(n23597), .CK(clk), .Q(n17217), .QN(n27296)
         );
  DFF_X2 avector23_reg_0__8_ ( .D(n23596), .CK(clk), .Q(n17254), .QN(n27295)
         );
  DFF_X2 avector23_reg_0__7_ ( .D(n23595), .CK(clk), .Q(n17291), .QN(n27294)
         );
  DFF_X2 avector23_reg_0__6_ ( .D(n23594), .CK(clk), .Q(n17328), .QN(n27293)
         );
  DFF_X2 avector23_reg_0__5_ ( .D(n23593), .CK(clk), .Q(n17365), .QN(n27292)
         );
  DFF_X2 avector23_reg_0__4_ ( .D(n23592), .CK(clk), .Q(n17402), .QN(n27291)
         );
  DFF_X2 avector23_reg_0__3_ ( .D(n23591), .CK(clk), .Q(n17439), .QN(n27290)
         );
  DFF_X2 avector23_reg_0__2_ ( .D(n23590), .CK(clk), .Q(n17476), .QN(n27289)
         );
  DFF_X2 avector23_reg_0__1_ ( .D(n23589), .CK(clk), .Q(n17513), .QN(n27288)
         );
  DFF_X2 avector23_reg_0__0_ ( .D(n23588), .CK(clk), .Q(n17550), .QN(n27287)
         );
  DFF_X2 avector22_reg_7__15_ ( .D(n23875), .CK(clk), .Q(n16973), .QN(n27622)
         );
  DFF_X2 avector22_reg_7__14_ ( .D(n23874), .CK(clk), .Q(n17010), .QN(n27621)
         );
  DFF_X2 avector22_reg_7__13_ ( .D(n23873), .CK(clk), .Q(n17047), .QN(n27620)
         );
  DFF_X2 avector22_reg_7__12_ ( .D(n23872), .CK(clk), .Q(n17084), .QN(n27619)
         );
  DFF_X2 avector22_reg_7__11_ ( .D(n23871), .CK(clk), .Q(n17121), .QN(n27618)
         );
  DFF_X2 avector22_reg_7__10_ ( .D(n23870), .CK(clk), .Q(n17158), .QN(n27617)
         );
  DFF_X2 avector22_reg_7__9_ ( .D(n23869), .CK(clk), .Q(n17195), .QN(n27616)
         );
  DFF_X2 avector22_reg_7__8_ ( .D(n23868), .CK(clk), .Q(n17232), .QN(n27615)
         );
  DFF_X2 avector22_reg_7__7_ ( .D(n23867), .CK(clk), .Q(n17269), .QN(n27614)
         );
  DFF_X2 avector22_reg_7__6_ ( .D(n23866), .CK(clk), .Q(n17306), .QN(n27613)
         );
  DFF_X2 avector22_reg_7__5_ ( .D(n23865), .CK(clk), .Q(n17343), .QN(n27612)
         );
  DFF_X2 avector22_reg_7__4_ ( .D(n23864), .CK(clk), .Q(n17380), .QN(n27611)
         );
  DFF_X2 avector22_reg_7__3_ ( .D(n23863), .CK(clk), .Q(n17417), .QN(n27610)
         );
  DFF_X2 avector22_reg_7__2_ ( .D(n23862), .CK(clk), .Q(n17454), .QN(n27609)
         );
  DFF_X2 avector22_reg_7__1_ ( .D(n23861), .CK(clk), .Q(n17491), .QN(n27608)
         );
  DFF_X2 avector22_reg_7__0_ ( .D(n23860), .CK(clk), .Q(n17528), .QN(n27607)
         );
  DFF_X2 avector22_reg_6__15_ ( .D(n23891), .CK(clk), .Q(n16971), .QN(n26854)
         );
  DFF_X2 avector22_reg_6__14_ ( .D(n23890), .CK(clk), .Q(n17008), .QN(n26853)
         );
  DFF_X2 avector22_reg_6__13_ ( .D(n23889), .CK(clk), .Q(n17045), .QN(n26852)
         );
  DFF_X2 avector22_reg_6__12_ ( .D(n23888), .CK(clk), .Q(n17082), .QN(n26851)
         );
  DFF_X2 avector22_reg_6__11_ ( .D(n23887), .CK(clk), .Q(n17119), .QN(n26850)
         );
  DFF_X2 avector22_reg_6__10_ ( .D(n23886), .CK(clk), .Q(n17156), .QN(n26849)
         );
  DFF_X2 avector22_reg_6__9_ ( .D(n23885), .CK(clk), .Q(n17193), .QN(n26848)
         );
  DFF_X2 avector22_reg_6__8_ ( .D(n23884), .CK(clk), .Q(n17230), .QN(n26847)
         );
  DFF_X2 avector22_reg_6__7_ ( .D(n23883), .CK(clk), .Q(n17267), .QN(n26846)
         );
  DFF_X2 avector22_reg_6__6_ ( .D(n23882), .CK(clk), .Q(n17304), .QN(n26845)
         );
  DFF_X2 avector22_reg_6__5_ ( .D(n23881), .CK(clk), .Q(n17341), .QN(n26844)
         );
  DFF_X2 avector22_reg_6__4_ ( .D(n23880), .CK(clk), .Q(n17378), .QN(n26843)
         );
  DFF_X2 avector22_reg_6__3_ ( .D(n23879), .CK(clk), .Q(n17415), .QN(n26842)
         );
  DFF_X2 avector22_reg_6__2_ ( .D(n23878), .CK(clk), .Q(n17452), .QN(n26841)
         );
  DFF_X2 avector22_reg_6__1_ ( .D(n23877), .CK(clk), .Q(n17489), .QN(n26840)
         );
  DFF_X2 avector22_reg_6__0_ ( .D(n23876), .CK(clk), .Q(n17526), .QN(n26839)
         );
  DFF_X2 avector22_reg_1__15_ ( .D(n23907), .CK(clk), .QN(n27110) );
  DFF_X2 avector22_reg_1__14_ ( .D(n23906), .CK(clk), .QN(n27109) );
  DFF_X2 avector22_reg_1__13_ ( .D(n23905), .CK(clk), .QN(n27108) );
  DFF_X2 avector22_reg_1__12_ ( .D(n23904), .CK(clk), .QN(n27107) );
  DFF_X2 avector22_reg_1__11_ ( .D(n23903), .CK(clk), .QN(n27106) );
  DFF_X2 avector22_reg_1__10_ ( .D(n23902), .CK(clk), .QN(n27105) );
  DFF_X2 avector22_reg_1__9_ ( .D(n23901), .CK(clk), .QN(n27104) );
  DFF_X2 avector22_reg_1__8_ ( .D(n23900), .CK(clk), .QN(n27103) );
  DFF_X2 avector22_reg_1__7_ ( .D(n23899), .CK(clk), .QN(n27102) );
  DFF_X2 avector22_reg_1__6_ ( .D(n23898), .CK(clk), .QN(n27101) );
  DFF_X2 avector22_reg_1__5_ ( .D(n23897), .CK(clk), .QN(n27100) );
  DFF_X2 avector22_reg_1__4_ ( .D(n23896), .CK(clk), .QN(n27099) );
  DFF_X2 avector22_reg_1__3_ ( .D(n23895), .CK(clk), .QN(n27098) );
  DFF_X2 avector22_reg_1__2_ ( .D(n23894), .CK(clk), .QN(n27097) );
  DFF_X2 avector22_reg_1__1_ ( .D(n23893), .CK(clk), .QN(n27096) );
  DFF_X2 avector22_reg_1__0_ ( .D(n23892), .CK(clk), .QN(n27095) );
  DFF_X2 avector22_reg_0__15_ ( .D(n23923), .CK(clk), .QN(n27366) );
  DFF_X2 avector22_reg_0__14_ ( .D(n23922), .CK(clk), .QN(n27365) );
  DFF_X2 avector22_reg_0__13_ ( .D(n23921), .CK(clk), .QN(n27364) );
  DFF_X2 avector22_reg_0__12_ ( .D(n23920), .CK(clk), .QN(n27363) );
  DFF_X2 avector22_reg_0__11_ ( .D(n23919), .CK(clk), .QN(n27362) );
  DFF_X2 avector22_reg_0__10_ ( .D(n23918), .CK(clk), .QN(n27361) );
  DFF_X2 avector22_reg_0__9_ ( .D(n23917), .CK(clk), .QN(n27360) );
  DFF_X2 avector22_reg_0__8_ ( .D(n23916), .CK(clk), .QN(n27359) );
  DFF_X2 avector22_reg_0__7_ ( .D(n23915), .CK(clk), .QN(n27358) );
  DFF_X2 avector22_reg_0__6_ ( .D(n23914), .CK(clk), .QN(n27357) );
  DFF_X2 avector22_reg_0__5_ ( .D(n23913), .CK(clk), .QN(n27356) );
  DFF_X2 avector22_reg_0__4_ ( .D(n23912), .CK(clk), .QN(n27355) );
  DFF_X2 avector22_reg_0__3_ ( .D(n23911), .CK(clk), .QN(n27354) );
  DFF_X2 avector22_reg_0__2_ ( .D(n23910), .CK(clk), .QN(n27353) );
  DFF_X2 avector22_reg_0__1_ ( .D(n23909), .CK(clk), .QN(n27352) );
  DFF_X2 avector22_reg_0__0_ ( .D(n23908), .CK(clk), .QN(n27351) );
  DFF_X2 avector21_reg_7__15_ ( .D(n24195), .CK(clk), .Q(n16982), .QN(n27686)
         );
  DFF_X2 avector21_reg_7__14_ ( .D(n24194), .CK(clk), .Q(n17019), .QN(n27685)
         );
  DFF_X2 avector21_reg_7__13_ ( .D(n24193), .CK(clk), .Q(n17056), .QN(n27684)
         );
  DFF_X2 avector21_reg_7__12_ ( .D(n24192), .CK(clk), .Q(n17093), .QN(n27683)
         );
  DFF_X2 avector21_reg_7__11_ ( .D(n24191), .CK(clk), .Q(n17130), .QN(n27682)
         );
  DFF_X2 avector21_reg_7__10_ ( .D(n24190), .CK(clk), .Q(n17167), .QN(n27681)
         );
  DFF_X2 avector21_reg_7__9_ ( .D(n24189), .CK(clk), .Q(n17204), .QN(n27680)
         );
  DFF_X2 avector21_reg_7__8_ ( .D(n24188), .CK(clk), .Q(n17241), .QN(n27679)
         );
  DFF_X2 avector21_reg_7__7_ ( .D(n24187), .CK(clk), .Q(n17278), .QN(n27678)
         );
  DFF_X2 avector21_reg_7__6_ ( .D(n24186), .CK(clk), .Q(n17315), .QN(n27677)
         );
  DFF_X2 avector21_reg_7__5_ ( .D(n24185), .CK(clk), .Q(n17352), .QN(n27676)
         );
  DFF_X2 avector21_reg_7__4_ ( .D(n24184), .CK(clk), .Q(n17389), .QN(n27675)
         );
  DFF_X2 avector21_reg_7__3_ ( .D(n24183), .CK(clk), .Q(n17426), .QN(n27674)
         );
  DFF_X2 avector21_reg_7__2_ ( .D(n24182), .CK(clk), .Q(n17463), .QN(n27673)
         );
  DFF_X2 avector21_reg_7__1_ ( .D(n24181), .CK(clk), .Q(n17500), .QN(n27672)
         );
  DFF_X2 avector21_reg_7__0_ ( .D(n24180), .CK(clk), .Q(n17537), .QN(n27671)
         );
  DFF_X2 avector21_reg_6__15_ ( .D(n24211), .CK(clk), .QN(n26918) );
  DFF_X2 avector21_reg_6__14_ ( .D(n24210), .CK(clk), .QN(n26917) );
  DFF_X2 avector21_reg_6__13_ ( .D(n24209), .CK(clk), .QN(n26916) );
  DFF_X2 avector21_reg_6__12_ ( .D(n24208), .CK(clk), .QN(n26915) );
  DFF_X2 avector21_reg_6__11_ ( .D(n24207), .CK(clk), .QN(n26914) );
  DFF_X2 avector21_reg_6__10_ ( .D(n24206), .CK(clk), .QN(n26913) );
  DFF_X2 avector21_reg_6__9_ ( .D(n24205), .CK(clk), .QN(n26912) );
  DFF_X2 avector21_reg_6__8_ ( .D(n24204), .CK(clk), .QN(n26911) );
  DFF_X2 avector21_reg_6__7_ ( .D(n24203), .CK(clk), .QN(n26910) );
  DFF_X2 avector21_reg_6__6_ ( .D(n24202), .CK(clk), .QN(n26909) );
  DFF_X2 avector21_reg_6__5_ ( .D(n24201), .CK(clk), .QN(n26908) );
  DFF_X2 avector21_reg_6__4_ ( .D(n24200), .CK(clk), .QN(n26907) );
  DFF_X2 avector21_reg_6__3_ ( .D(n24199), .CK(clk), .QN(n26906) );
  DFF_X2 avector21_reg_6__2_ ( .D(n24198), .CK(clk), .QN(n26905) );
  DFF_X2 avector21_reg_6__1_ ( .D(n24197), .CK(clk), .QN(n26904) );
  DFF_X2 avector21_reg_6__0_ ( .D(n24196), .CK(clk), .QN(n26903) );
  DFF_X2 avector21_reg_1__15_ ( .D(n24227), .CK(clk), .QN(n27174) );
  DFF_X2 avector21_reg_1__14_ ( .D(n24226), .CK(clk), .QN(n27173) );
  DFF_X2 avector21_reg_1__13_ ( .D(n24225), .CK(clk), .QN(n27172) );
  DFF_X2 avector21_reg_1__12_ ( .D(n24224), .CK(clk), .QN(n27171) );
  DFF_X2 avector21_reg_1__11_ ( .D(n24223), .CK(clk), .QN(n27170) );
  DFF_X2 avector21_reg_1__10_ ( .D(n24222), .CK(clk), .QN(n27169) );
  DFF_X2 avector21_reg_1__9_ ( .D(n24221), .CK(clk), .QN(n27168) );
  DFF_X2 avector21_reg_1__8_ ( .D(n24220), .CK(clk), .QN(n27167) );
  DFF_X2 avector21_reg_1__7_ ( .D(n24219), .CK(clk), .QN(n27166) );
  DFF_X2 avector21_reg_1__6_ ( .D(n24218), .CK(clk), .QN(n27165) );
  DFF_X2 avector21_reg_1__5_ ( .D(n24217), .CK(clk), .QN(n27164) );
  DFF_X2 avector21_reg_1__4_ ( .D(n24216), .CK(clk), .QN(n27163) );
  DFF_X2 avector21_reg_1__3_ ( .D(n24215), .CK(clk), .QN(n27162) );
  DFF_X2 avector21_reg_1__2_ ( .D(n24214), .CK(clk), .QN(n27161) );
  DFF_X2 avector21_reg_1__1_ ( .D(n24213), .CK(clk), .QN(n27160) );
  DFF_X2 avector21_reg_1__0_ ( .D(n24212), .CK(clk), .QN(n27159) );
  DFF_X2 avector21_reg_0__15_ ( .D(n24243), .CK(clk), .QN(n27430) );
  DFF_X2 avector21_reg_0__14_ ( .D(n24242), .CK(clk), .QN(n27429) );
  DFF_X2 avector21_reg_0__13_ ( .D(n24241), .CK(clk), .QN(n27428) );
  DFF_X2 avector21_reg_0__12_ ( .D(n24240), .CK(clk), .QN(n27427) );
  DFF_X2 avector21_reg_0__11_ ( .D(n24239), .CK(clk), .QN(n27426) );
  DFF_X2 avector21_reg_0__10_ ( .D(n24238), .CK(clk), .QN(n27425) );
  DFF_X2 avector21_reg_0__9_ ( .D(n24237), .CK(clk), .QN(n27424) );
  DFF_X2 avector21_reg_0__8_ ( .D(n24236), .CK(clk), .QN(n27423) );
  DFF_X2 avector21_reg_0__7_ ( .D(n24235), .CK(clk), .QN(n27422) );
  DFF_X2 avector21_reg_0__6_ ( .D(n24234), .CK(clk), .QN(n27421) );
  DFF_X2 avector21_reg_0__5_ ( .D(n24233), .CK(clk), .QN(n27420) );
  DFF_X2 avector21_reg_0__4_ ( .D(n24232), .CK(clk), .QN(n27419) );
  DFF_X2 avector21_reg_0__3_ ( .D(n24231), .CK(clk), .QN(n27418) );
  DFF_X2 avector21_reg_0__2_ ( .D(n24230), .CK(clk), .QN(n27417) );
  DFF_X2 avector21_reg_0__1_ ( .D(n24229), .CK(clk), .QN(n27416) );
  DFF_X2 avector21_reg_0__0_ ( .D(n24228), .CK(clk), .QN(n27415) );
  DFF_X2 avector20_reg_7__15_ ( .D(n24515), .CK(clk), .QN(n27750) );
  DFF_X2 avector20_reg_7__14_ ( .D(n24514), .CK(clk), .QN(n27749) );
  DFF_X2 avector20_reg_7__13_ ( .D(n24513), .CK(clk), .QN(n27748) );
  DFF_X2 avector20_reg_7__12_ ( .D(n24512), .CK(clk), .QN(n27747) );
  DFF_X2 avector20_reg_7__11_ ( .D(n24511), .CK(clk), .QN(n27746) );
  DFF_X2 avector20_reg_7__10_ ( .D(n24510), .CK(clk), .QN(n27745) );
  DFF_X2 avector20_reg_7__9_ ( .D(n24509), .CK(clk), .QN(n27744) );
  DFF_X2 avector20_reg_7__8_ ( .D(n24508), .CK(clk), .QN(n27743) );
  DFF_X2 avector20_reg_7__7_ ( .D(n24507), .CK(clk), .QN(n27742) );
  DFF_X2 avector20_reg_7__6_ ( .D(n24506), .CK(clk), .QN(n27741) );
  DFF_X2 avector20_reg_7__5_ ( .D(n24505), .CK(clk), .QN(n27740) );
  DFF_X2 avector20_reg_7__4_ ( .D(n24504), .CK(clk), .QN(n27739) );
  DFF_X2 avector20_reg_7__3_ ( .D(n24503), .CK(clk), .QN(n27738) );
  DFF_X2 avector20_reg_7__2_ ( .D(n24502), .CK(clk), .QN(n27737) );
  DFF_X2 avector20_reg_7__1_ ( .D(n24501), .CK(clk), .QN(n27736) );
  DFF_X2 avector20_reg_7__0_ ( .D(n24500), .CK(clk), .QN(n27735) );
  DFF_X2 avector20_reg_6__15_ ( .D(n24531), .CK(clk), .QN(n26982) );
  DFF_X2 avector20_reg_6__14_ ( .D(n24530), .CK(clk), .QN(n26981) );
  DFF_X2 avector20_reg_6__13_ ( .D(n24529), .CK(clk), .QN(n26980) );
  DFF_X2 avector20_reg_6__12_ ( .D(n24528), .CK(clk), .QN(n26979) );
  DFF_X2 avector20_reg_6__11_ ( .D(n24527), .CK(clk), .QN(n26978) );
  DFF_X2 avector20_reg_6__10_ ( .D(n24526), .CK(clk), .QN(n26977) );
  DFF_X2 avector20_reg_6__9_ ( .D(n24525), .CK(clk), .QN(n26976) );
  DFF_X2 avector20_reg_6__8_ ( .D(n24524), .CK(clk), .QN(n26975) );
  DFF_X2 avector20_reg_6__7_ ( .D(n24523), .CK(clk), .QN(n26974) );
  DFF_X2 avector20_reg_6__6_ ( .D(n24522), .CK(clk), .QN(n26973) );
  DFF_X2 avector20_reg_6__5_ ( .D(n24521), .CK(clk), .QN(n26972) );
  DFF_X2 avector20_reg_6__4_ ( .D(n24520), .CK(clk), .QN(n26971) );
  DFF_X2 avector20_reg_6__3_ ( .D(n24519), .CK(clk), .QN(n26970) );
  DFF_X2 avector20_reg_6__2_ ( .D(n24518), .CK(clk), .QN(n26969) );
  DFF_X2 avector20_reg_6__1_ ( .D(n24517), .CK(clk), .QN(n26968) );
  DFF_X2 avector20_reg_6__0_ ( .D(n24516), .CK(clk), .QN(n26967) );
  DFF_X2 avector20_reg_1__15_ ( .D(n24547), .CK(clk), .Q(n16985), .QN(n27238)
         );
  DFF_X2 avector20_reg_1__14_ ( .D(n24546), .CK(clk), .Q(n17022), .QN(n27237)
         );
  DFF_X2 avector20_reg_1__13_ ( .D(n24545), .CK(clk), .Q(n17059), .QN(n27236)
         );
  DFF_X2 avector20_reg_1__12_ ( .D(n24544), .CK(clk), .Q(n17096), .QN(n27235)
         );
  DFF_X2 avector20_reg_1__11_ ( .D(n24543), .CK(clk), .Q(n17133), .QN(n27234)
         );
  DFF_X2 avector20_reg_1__10_ ( .D(n24542), .CK(clk), .Q(n17170), .QN(n27233)
         );
  DFF_X2 avector20_reg_1__9_ ( .D(n24541), .CK(clk), .Q(n17207), .QN(n27232)
         );
  DFF_X2 avector20_reg_1__8_ ( .D(n24540), .CK(clk), .Q(n17244), .QN(n27231)
         );
  DFF_X2 avector20_reg_1__7_ ( .D(n24539), .CK(clk), .Q(n17281), .QN(n27230)
         );
  DFF_X2 avector20_reg_1__6_ ( .D(n24538), .CK(clk), .Q(n17318), .QN(n27229)
         );
  DFF_X2 avector20_reg_1__5_ ( .D(n24537), .CK(clk), .Q(n17355), .QN(n27228)
         );
  DFF_X2 avector20_reg_1__4_ ( .D(n24536), .CK(clk), .Q(n17392), .QN(n27227)
         );
  DFF_X2 avector20_reg_1__3_ ( .D(n24535), .CK(clk), .Q(n17429), .QN(n27226)
         );
  DFF_X2 avector20_reg_1__2_ ( .D(n24534), .CK(clk), .Q(n17466), .QN(n27225)
         );
  DFF_X2 avector20_reg_1__1_ ( .D(n24533), .CK(clk), .Q(n17503), .QN(n27224)
         );
  DFF_X2 avector20_reg_1__0_ ( .D(n24532), .CK(clk), .Q(n17540), .QN(n27223)
         );
  DFF_X2 avector20_reg_0__15_ ( .D(n24563), .CK(clk), .Q(n16986), .QN(n27494)
         );
  DFF_X2 avector20_reg_0__14_ ( .D(n24562), .CK(clk), .Q(n17023), .QN(n27493)
         );
  DFF_X2 avector20_reg_0__13_ ( .D(n24561), .CK(clk), .Q(n17060), .QN(n27492)
         );
  DFF_X2 avector20_reg_0__12_ ( .D(n24560), .CK(clk), .Q(n17097), .QN(n27491)
         );
  DFF_X2 avector20_reg_0__11_ ( .D(n24559), .CK(clk), .Q(n17134), .QN(n27490)
         );
  DFF_X2 avector20_reg_0__10_ ( .D(n24558), .CK(clk), .Q(n17171), .QN(n27489)
         );
  DFF_X2 avector20_reg_0__9_ ( .D(n24557), .CK(clk), .Q(n17208), .QN(n27488)
         );
  DFF_X2 avector20_reg_0__8_ ( .D(n24556), .CK(clk), .Q(n17245), .QN(n27487)
         );
  DFF_X2 avector20_reg_0__7_ ( .D(n24555), .CK(clk), .Q(n17282), .QN(n27486)
         );
  DFF_X2 avector20_reg_0__6_ ( .D(n24554), .CK(clk), .Q(n17319), .QN(n27485)
         );
  DFF_X2 avector20_reg_0__5_ ( .D(n24553), .CK(clk), .Q(n17356), .QN(n27484)
         );
  DFF_X2 avector20_reg_0__4_ ( .D(n24552), .CK(clk), .Q(n17393), .QN(n27483)
         );
  DFF_X2 avector20_reg_0__3_ ( .D(n24551), .CK(clk), .Q(n17430), .QN(n27482)
         );
  DFF_X2 avector20_reg_0__2_ ( .D(n24550), .CK(clk), .Q(n17467), .QN(n27481)
         );
  DFF_X2 avector20_reg_0__1_ ( .D(n24549), .CK(clk), .Q(n17504), .QN(n27480)
         );
  DFF_X2 avector20_reg_0__0_ ( .D(n24548), .CK(clk), .Q(n17541), .QN(n27479)
         );
  DFF_X2 avector13_reg_7__15_ ( .D(n23635), .CK(clk), .QN(n27574) );
  DFF_X2 avector13_reg_7__14_ ( .D(n23634), .CK(clk), .QN(n27573) );
  DFF_X2 avector13_reg_7__13_ ( .D(n23633), .CK(clk), .QN(n27572) );
  DFF_X2 avector13_reg_7__12_ ( .D(n23632), .CK(clk), .QN(n27571) );
  DFF_X2 avector13_reg_7__11_ ( .D(n23631), .CK(clk), .QN(n27570) );
  DFF_X2 avector13_reg_7__10_ ( .D(n23630), .CK(clk), .QN(n27569) );
  DFF_X2 avector13_reg_7__9_ ( .D(n23629), .CK(clk), .QN(n27568) );
  DFF_X2 avector13_reg_7__8_ ( .D(n23628), .CK(clk), .QN(n27567) );
  DFF_X2 avector13_reg_7__7_ ( .D(n23627), .CK(clk), .QN(n27566) );
  DFF_X2 avector13_reg_7__6_ ( .D(n23626), .CK(clk), .QN(n27565) );
  DFF_X2 avector13_reg_7__5_ ( .D(n23625), .CK(clk), .QN(n27564) );
  DFF_X2 avector13_reg_7__4_ ( .D(n23624), .CK(clk), .QN(n27563) );
  DFF_X2 avector13_reg_7__3_ ( .D(n23623), .CK(clk), .QN(n27562) );
  DFF_X2 avector13_reg_7__2_ ( .D(n23622), .CK(clk), .QN(n27561) );
  DFF_X2 avector13_reg_7__1_ ( .D(n23621), .CK(clk), .QN(n27560) );
  DFF_X2 avector13_reg_7__0_ ( .D(n23620), .CK(clk), .QN(n27559) );
  DFF_X2 avector13_reg_6__15_ ( .D(n23651), .CK(clk), .QN(n26806) );
  DFF_X2 avector13_reg_6__14_ ( .D(n23650), .CK(clk), .QN(n26805) );
  DFF_X2 avector13_reg_6__13_ ( .D(n23649), .CK(clk), .QN(n26804) );
  DFF_X2 avector13_reg_6__12_ ( .D(n23648), .CK(clk), .QN(n26803) );
  DFF_X2 avector13_reg_6__11_ ( .D(n23647), .CK(clk), .QN(n26802) );
  DFF_X2 avector13_reg_6__10_ ( .D(n23646), .CK(clk), .QN(n26801) );
  DFF_X2 avector13_reg_6__9_ ( .D(n23645), .CK(clk), .QN(n26800) );
  DFF_X2 avector13_reg_6__8_ ( .D(n23644), .CK(clk), .QN(n26799) );
  DFF_X2 avector13_reg_6__7_ ( .D(n23643), .CK(clk), .QN(n26798) );
  DFF_X2 avector13_reg_6__6_ ( .D(n23642), .CK(clk), .QN(n26797) );
  DFF_X2 avector13_reg_6__5_ ( .D(n23641), .CK(clk), .QN(n26796) );
  DFF_X2 avector13_reg_6__4_ ( .D(n23640), .CK(clk), .QN(n26795) );
  DFF_X2 avector13_reg_6__3_ ( .D(n23639), .CK(clk), .QN(n26794) );
  DFF_X2 avector13_reg_6__2_ ( .D(n23638), .CK(clk), .QN(n26793) );
  DFF_X2 avector13_reg_6__1_ ( .D(n23637), .CK(clk), .QN(n26792) );
  DFF_X2 avector13_reg_6__0_ ( .D(n23636), .CK(clk), .QN(n26791) );
  DFF_X2 avector13_reg_1__15_ ( .D(n23667), .CK(clk), .Q(n17586), .QN(n27062)
         );
  DFF_X2 avector13_reg_1__14_ ( .D(n23666), .CK(clk), .Q(n17623), .QN(n27061)
         );
  DFF_X2 avector13_reg_1__13_ ( .D(n23665), .CK(clk), .Q(n17660), .QN(n27060)
         );
  DFF_X2 avector13_reg_1__12_ ( .D(n23664), .CK(clk), .Q(n17697), .QN(n27059)
         );
  DFF_X2 avector13_reg_1__11_ ( .D(n23663), .CK(clk), .Q(n17734), .QN(n27058)
         );
  DFF_X2 avector13_reg_1__10_ ( .D(n23662), .CK(clk), .Q(n17771), .QN(n27057)
         );
  DFF_X2 avector13_reg_1__9_ ( .D(n23661), .CK(clk), .Q(n17808), .QN(n27056)
         );
  DFF_X2 avector13_reg_1__8_ ( .D(n23660), .CK(clk), .Q(n17845), .QN(n27055)
         );
  DFF_X2 avector13_reg_1__7_ ( .D(n23659), .CK(clk), .Q(n17882), .QN(n27054)
         );
  DFF_X2 avector13_reg_1__6_ ( .D(n23658), .CK(clk), .Q(n17919), .QN(n27053)
         );
  DFF_X2 avector13_reg_1__5_ ( .D(n23657), .CK(clk), .Q(n17956), .QN(n27052)
         );
  DFF_X2 avector13_reg_1__4_ ( .D(n23656), .CK(clk), .Q(n17993), .QN(n27051)
         );
  DFF_X2 avector13_reg_1__3_ ( .D(n23655), .CK(clk), .Q(n18030), .QN(n27050)
         );
  DFF_X2 avector13_reg_1__2_ ( .D(n23654), .CK(clk), .Q(n18067), .QN(n27049)
         );
  DFF_X2 avector13_reg_1__1_ ( .D(n23653), .CK(clk), .Q(n18104), .QN(n27048)
         );
  DFF_X2 avector13_reg_1__0_ ( .D(n23652), .CK(clk), .Q(n18141), .QN(n27047)
         );
  DFF_X2 avector13_reg_0__15_ ( .D(n23683), .CK(clk), .Q(n17587), .QN(n27318)
         );
  DFF_X2 avector13_reg_0__14_ ( .D(n23682), .CK(clk), .Q(n17624), .QN(n27317)
         );
  DFF_X2 avector13_reg_0__13_ ( .D(n23681), .CK(clk), .Q(n17661), .QN(n27316)
         );
  DFF_X2 avector13_reg_0__12_ ( .D(n23680), .CK(clk), .Q(n17698), .QN(n27315)
         );
  DFF_X2 avector13_reg_0__11_ ( .D(n23679), .CK(clk), .Q(n17735), .QN(n27314)
         );
  DFF_X2 avector13_reg_0__10_ ( .D(n23678), .CK(clk), .Q(n17772), .QN(n27313)
         );
  DFF_X2 avector13_reg_0__9_ ( .D(n23677), .CK(clk), .Q(n17809), .QN(n27312)
         );
  DFF_X2 avector13_reg_0__8_ ( .D(n23676), .CK(clk), .Q(n17846), .QN(n27311)
         );
  DFF_X2 avector13_reg_0__7_ ( .D(n23675), .CK(clk), .Q(n17883), .QN(n27310)
         );
  DFF_X2 avector13_reg_0__6_ ( .D(n23674), .CK(clk), .Q(n17920), .QN(n27309)
         );
  DFF_X2 avector13_reg_0__5_ ( .D(n23673), .CK(clk), .Q(n17957), .QN(n27308)
         );
  DFF_X2 avector13_reg_0__4_ ( .D(n23672), .CK(clk), .Q(n17994), .QN(n27307)
         );
  DFF_X2 avector13_reg_0__3_ ( .D(n23671), .CK(clk), .Q(n18031), .QN(n27306)
         );
  DFF_X2 avector13_reg_0__2_ ( .D(n23670), .CK(clk), .Q(n18068), .QN(n27305)
         );
  DFF_X2 avector13_reg_0__1_ ( .D(n23669), .CK(clk), .Q(n18105), .QN(n27304)
         );
  DFF_X2 avector13_reg_0__0_ ( .D(n23668), .CK(clk), .Q(n18142), .QN(n27303)
         );
  DFF_X2 avector12_reg_7__15_ ( .D(n23955), .CK(clk), .Q(n17565), .QN(n27638)
         );
  DFF_X2 avector12_reg_7__14_ ( .D(n23954), .CK(clk), .Q(n17602), .QN(n27637)
         );
  DFF_X2 avector12_reg_7__13_ ( .D(n23953), .CK(clk), .Q(n17639), .QN(n27636)
         );
  DFF_X2 avector12_reg_7__12_ ( .D(n23952), .CK(clk), .Q(n17676), .QN(n27635)
         );
  DFF_X2 avector12_reg_7__11_ ( .D(n23951), .CK(clk), .Q(n17713), .QN(n27634)
         );
  DFF_X2 avector12_reg_7__10_ ( .D(n23950), .CK(clk), .Q(n17750), .QN(n27633)
         );
  DFF_X2 avector12_reg_7__9_ ( .D(n23949), .CK(clk), .Q(n17787), .QN(n27632)
         );
  DFF_X2 avector12_reg_7__8_ ( .D(n23948), .CK(clk), .Q(n17824), .QN(n27631)
         );
  DFF_X2 avector12_reg_7__7_ ( .D(n23947), .CK(clk), .Q(n17861), .QN(n27630)
         );
  DFF_X2 avector12_reg_7__6_ ( .D(n23946), .CK(clk), .Q(n17898), .QN(n27629)
         );
  DFF_X2 avector12_reg_7__5_ ( .D(n23945), .CK(clk), .Q(n17935), .QN(n27628)
         );
  DFF_X2 avector12_reg_7__4_ ( .D(n23944), .CK(clk), .Q(n17972), .QN(n27627)
         );
  DFF_X2 avector12_reg_7__3_ ( .D(n23943), .CK(clk), .Q(n18009), .QN(n27626)
         );
  DFF_X2 avector12_reg_7__2_ ( .D(n23942), .CK(clk), .Q(n18046), .QN(n27625)
         );
  DFF_X2 avector12_reg_7__1_ ( .D(n23941), .CK(clk), .Q(n18083), .QN(n27624)
         );
  DFF_X2 avector12_reg_7__0_ ( .D(n23940), .CK(clk), .Q(n18120), .QN(n27623)
         );
  DFF_X2 avector12_reg_6__15_ ( .D(n23971), .CK(clk), .Q(n17563), .QN(n26870)
         );
  DFF_X2 avector12_reg_6__14_ ( .D(n23970), .CK(clk), .Q(n17600), .QN(n26869)
         );
  DFF_X2 avector12_reg_6__13_ ( .D(n23969), .CK(clk), .Q(n17637), .QN(n26868)
         );
  DFF_X2 avector12_reg_6__12_ ( .D(n23968), .CK(clk), .Q(n17674), .QN(n26867)
         );
  DFF_X2 avector12_reg_6__11_ ( .D(n23967), .CK(clk), .Q(n17711), .QN(n26866)
         );
  DFF_X2 avector12_reg_6__10_ ( .D(n23966), .CK(clk), .Q(n17748), .QN(n26865)
         );
  DFF_X2 avector12_reg_6__9_ ( .D(n23965), .CK(clk), .Q(n17785), .QN(n26864)
         );
  DFF_X2 avector12_reg_6__8_ ( .D(n23964), .CK(clk), .Q(n17822), .QN(n26863)
         );
  DFF_X2 avector12_reg_6__7_ ( .D(n23963), .CK(clk), .Q(n17859), .QN(n26862)
         );
  DFF_X2 avector12_reg_6__6_ ( .D(n23962), .CK(clk), .Q(n17896), .QN(n26861)
         );
  DFF_X2 avector12_reg_6__5_ ( .D(n23961), .CK(clk), .Q(n17933), .QN(n26860)
         );
  DFF_X2 avector12_reg_6__4_ ( .D(n23960), .CK(clk), .Q(n17970), .QN(n26859)
         );
  DFF_X2 avector12_reg_6__3_ ( .D(n23959), .CK(clk), .Q(n18007), .QN(n26858)
         );
  DFF_X2 avector12_reg_6__2_ ( .D(n23958), .CK(clk), .Q(n18044), .QN(n26857)
         );
  DFF_X2 avector12_reg_6__1_ ( .D(n23957), .CK(clk), .Q(n18081), .QN(n26856)
         );
  DFF_X2 avector12_reg_6__0_ ( .D(n23956), .CK(clk), .Q(n18118), .QN(n26855)
         );
  DFF_X2 avector12_reg_1__15_ ( .D(n23987), .CK(clk), .QN(n27126) );
  DFF_X2 avector12_reg_1__14_ ( .D(n23986), .CK(clk), .QN(n27125) );
  DFF_X2 avector12_reg_1__13_ ( .D(n23985), .CK(clk), .QN(n27124) );
  DFF_X2 avector12_reg_1__12_ ( .D(n23984), .CK(clk), .QN(n27123) );
  DFF_X2 avector12_reg_1__11_ ( .D(n23983), .CK(clk), .QN(n27122) );
  DFF_X2 avector12_reg_1__10_ ( .D(n23982), .CK(clk), .QN(n27121) );
  DFF_X2 avector12_reg_1__9_ ( .D(n23981), .CK(clk), .QN(n27120) );
  DFF_X2 avector12_reg_1__8_ ( .D(n23980), .CK(clk), .QN(n27119) );
  DFF_X2 avector12_reg_1__7_ ( .D(n23979), .CK(clk), .QN(n27118) );
  DFF_X2 avector12_reg_1__6_ ( .D(n23978), .CK(clk), .QN(n27117) );
  DFF_X2 avector12_reg_1__5_ ( .D(n23977), .CK(clk), .QN(n27116) );
  DFF_X2 avector12_reg_1__4_ ( .D(n23976), .CK(clk), .QN(n27115) );
  DFF_X2 avector12_reg_1__3_ ( .D(n23975), .CK(clk), .QN(n27114) );
  DFF_X2 avector12_reg_1__2_ ( .D(n23974), .CK(clk), .QN(n27113) );
  DFF_X2 avector12_reg_1__1_ ( .D(n23973), .CK(clk), .QN(n27112) );
  DFF_X2 avector12_reg_1__0_ ( .D(n23972), .CK(clk), .QN(n27111) );
  DFF_X2 avector12_reg_0__15_ ( .D(n24003), .CK(clk), .QN(n27382) );
  DFF_X2 avector12_reg_0__14_ ( .D(n24002), .CK(clk), .QN(n27381) );
  DFF_X2 avector12_reg_0__13_ ( .D(n24001), .CK(clk), .QN(n27380) );
  DFF_X2 avector12_reg_0__12_ ( .D(n24000), .CK(clk), .QN(n27379) );
  DFF_X2 avector12_reg_0__11_ ( .D(n23999), .CK(clk), .QN(n27378) );
  DFF_X2 avector12_reg_0__10_ ( .D(n23998), .CK(clk), .QN(n27377) );
  DFF_X2 avector12_reg_0__9_ ( .D(n23997), .CK(clk), .QN(n27376) );
  DFF_X2 avector12_reg_0__8_ ( .D(n23996), .CK(clk), .QN(n27375) );
  DFF_X2 avector12_reg_0__7_ ( .D(n23995), .CK(clk), .QN(n27374) );
  DFF_X2 avector12_reg_0__6_ ( .D(n23994), .CK(clk), .QN(n27373) );
  DFF_X2 avector12_reg_0__5_ ( .D(n23993), .CK(clk), .QN(n27372) );
  DFF_X2 avector12_reg_0__4_ ( .D(n23992), .CK(clk), .QN(n27371) );
  DFF_X2 avector12_reg_0__3_ ( .D(n23991), .CK(clk), .QN(n27370) );
  DFF_X2 avector12_reg_0__2_ ( .D(n23990), .CK(clk), .QN(n27369) );
  DFF_X2 avector12_reg_0__1_ ( .D(n23989), .CK(clk), .QN(n27368) );
  DFF_X2 avector12_reg_0__0_ ( .D(n23988), .CK(clk), .QN(n27367) );
  DFF_X2 avector11_reg_7__15_ ( .D(n24275), .CK(clk), .Q(n17574), .QN(n27702)
         );
  DFF_X2 avector11_reg_7__14_ ( .D(n24274), .CK(clk), .Q(n17611), .QN(n27701)
         );
  DFF_X2 avector11_reg_7__13_ ( .D(n24273), .CK(clk), .Q(n17648), .QN(n27700)
         );
  DFF_X2 avector11_reg_7__12_ ( .D(n24272), .CK(clk), .Q(n17685), .QN(n27699)
         );
  DFF_X2 avector11_reg_7__11_ ( .D(n24271), .CK(clk), .Q(n17722), .QN(n27698)
         );
  DFF_X2 avector11_reg_7__10_ ( .D(n24270), .CK(clk), .Q(n17759), .QN(n27697)
         );
  DFF_X2 avector11_reg_7__9_ ( .D(n24269), .CK(clk), .Q(n17796), .QN(n27696)
         );
  DFF_X2 avector11_reg_7__8_ ( .D(n24268), .CK(clk), .Q(n17833), .QN(n27695)
         );
  DFF_X2 avector11_reg_7__7_ ( .D(n24267), .CK(clk), .Q(n17870), .QN(n27694)
         );
  DFF_X2 avector11_reg_7__6_ ( .D(n24266), .CK(clk), .Q(n17907), .QN(n27693)
         );
  DFF_X2 avector11_reg_7__5_ ( .D(n24265), .CK(clk), .Q(n17944), .QN(n27692)
         );
  DFF_X2 avector11_reg_7__4_ ( .D(n24264), .CK(clk), .Q(n17981), .QN(n27691)
         );
  DFF_X2 avector11_reg_7__3_ ( .D(n24263), .CK(clk), .Q(n18018), .QN(n27690)
         );
  DFF_X2 avector11_reg_7__2_ ( .D(n24262), .CK(clk), .Q(n18055), .QN(n27689)
         );
  DFF_X2 avector11_reg_7__1_ ( .D(n24261), .CK(clk), .Q(n18092), .QN(n27688)
         );
  DFF_X2 avector11_reg_7__0_ ( .D(n24260), .CK(clk), .Q(n18129), .QN(n27687)
         );
  DFF_X2 avector11_reg_6__15_ ( .D(n24291), .CK(clk), .QN(n26934) );
  DFF_X2 avector11_reg_6__14_ ( .D(n24290), .CK(clk), .QN(n26933) );
  DFF_X2 avector11_reg_6__13_ ( .D(n24289), .CK(clk), .QN(n26932) );
  DFF_X2 avector11_reg_6__12_ ( .D(n24288), .CK(clk), .QN(n26931) );
  DFF_X2 avector11_reg_6__11_ ( .D(n24287), .CK(clk), .QN(n26930) );
  DFF_X2 avector11_reg_6__10_ ( .D(n24286), .CK(clk), .QN(n26929) );
  DFF_X2 avector11_reg_6__9_ ( .D(n24285), .CK(clk), .QN(n26928) );
  DFF_X2 avector11_reg_6__8_ ( .D(n24284), .CK(clk), .QN(n26927) );
  DFF_X2 avector11_reg_6__7_ ( .D(n24283), .CK(clk), .QN(n26926) );
  DFF_X2 avector11_reg_6__6_ ( .D(n24282), .CK(clk), .QN(n26925) );
  DFF_X2 avector11_reg_6__5_ ( .D(n24281), .CK(clk), .QN(n26924) );
  DFF_X2 avector11_reg_6__4_ ( .D(n24280), .CK(clk), .QN(n26923) );
  DFF_X2 avector11_reg_6__3_ ( .D(n24279), .CK(clk), .QN(n26922) );
  DFF_X2 avector11_reg_6__2_ ( .D(n24278), .CK(clk), .QN(n26921) );
  DFF_X2 avector11_reg_6__1_ ( .D(n24277), .CK(clk), .QN(n26920) );
  DFF_X2 avector11_reg_6__0_ ( .D(n24276), .CK(clk), .QN(n26919) );
  DFF_X2 avector11_reg_1__15_ ( .D(n24307), .CK(clk), .QN(n27190) );
  DFF_X2 avector11_reg_1__14_ ( .D(n24306), .CK(clk), .QN(n27189) );
  DFF_X2 avector11_reg_1__13_ ( .D(n24305), .CK(clk), .QN(n27188) );
  DFF_X2 avector11_reg_1__12_ ( .D(n24304), .CK(clk), .QN(n27187) );
  DFF_X2 avector11_reg_1__11_ ( .D(n24303), .CK(clk), .QN(n27186) );
  DFF_X2 avector11_reg_1__10_ ( .D(n24302), .CK(clk), .QN(n27185) );
  DFF_X2 avector11_reg_1__9_ ( .D(n24301), .CK(clk), .QN(n27184) );
  DFF_X2 avector11_reg_1__8_ ( .D(n24300), .CK(clk), .QN(n27183) );
  DFF_X2 avector11_reg_1__7_ ( .D(n24299), .CK(clk), .QN(n27182) );
  DFF_X2 avector11_reg_1__6_ ( .D(n24298), .CK(clk), .QN(n27181) );
  DFF_X2 avector11_reg_1__5_ ( .D(n24297), .CK(clk), .QN(n27180) );
  DFF_X2 avector11_reg_1__4_ ( .D(n24296), .CK(clk), .QN(n27179) );
  DFF_X2 avector11_reg_1__3_ ( .D(n24295), .CK(clk), .QN(n27178) );
  DFF_X2 avector11_reg_1__2_ ( .D(n24294), .CK(clk), .QN(n27177) );
  DFF_X2 avector11_reg_1__1_ ( .D(n24293), .CK(clk), .QN(n27176) );
  DFF_X2 avector11_reg_1__0_ ( .D(n24292), .CK(clk), .QN(n27175) );
  DFF_X2 avector11_reg_0__15_ ( .D(n24323), .CK(clk), .QN(n27446) );
  DFF_X2 avector11_reg_0__14_ ( .D(n24322), .CK(clk), .QN(n27445) );
  DFF_X2 avector11_reg_0__13_ ( .D(n24321), .CK(clk), .QN(n27444) );
  DFF_X2 avector11_reg_0__12_ ( .D(n24320), .CK(clk), .QN(n27443) );
  DFF_X2 avector11_reg_0__11_ ( .D(n24319), .CK(clk), .QN(n27442) );
  DFF_X2 avector11_reg_0__10_ ( .D(n24318), .CK(clk), .QN(n27441) );
  DFF_X2 avector11_reg_0__9_ ( .D(n24317), .CK(clk), .QN(n27440) );
  DFF_X2 avector11_reg_0__8_ ( .D(n24316), .CK(clk), .QN(n27439) );
  DFF_X2 avector11_reg_0__7_ ( .D(n24315), .CK(clk), .QN(n27438) );
  DFF_X2 avector11_reg_0__6_ ( .D(n24314), .CK(clk), .QN(n27437) );
  DFF_X2 avector11_reg_0__5_ ( .D(n24313), .CK(clk), .QN(n27436) );
  DFF_X2 avector11_reg_0__4_ ( .D(n24312), .CK(clk), .QN(n27435) );
  DFF_X2 avector11_reg_0__3_ ( .D(n24311), .CK(clk), .QN(n27434) );
  DFF_X2 avector11_reg_0__2_ ( .D(n24310), .CK(clk), .QN(n27433) );
  DFF_X2 avector11_reg_0__1_ ( .D(n24309), .CK(clk), .QN(n27432) );
  DFF_X2 avector11_reg_0__0_ ( .D(n24308), .CK(clk), .QN(n27431) );
  DFF_X2 avector10_reg_7__15_ ( .D(n24595), .CK(clk), .QN(n27766) );
  DFF_X2 avector10_reg_7__14_ ( .D(n24594), .CK(clk), .QN(n27765) );
  DFF_X2 avector10_reg_7__13_ ( .D(n24593), .CK(clk), .QN(n27764) );
  DFF_X2 avector10_reg_7__12_ ( .D(n24592), .CK(clk), .QN(n27763) );
  DFF_X2 avector10_reg_7__11_ ( .D(n24591), .CK(clk), .QN(n27762) );
  DFF_X2 avector10_reg_7__10_ ( .D(n24590), .CK(clk), .QN(n27761) );
  DFF_X2 avector10_reg_7__9_ ( .D(n24589), .CK(clk), .QN(n27760) );
  DFF_X2 avector10_reg_7__8_ ( .D(n24588), .CK(clk), .QN(n27759) );
  DFF_X2 avector10_reg_7__7_ ( .D(n24587), .CK(clk), .QN(n27758) );
  DFF_X2 avector10_reg_7__6_ ( .D(n24586), .CK(clk), .QN(n27757) );
  DFF_X2 avector10_reg_7__5_ ( .D(n24585), .CK(clk), .QN(n27756) );
  DFF_X2 avector10_reg_7__4_ ( .D(n24584), .CK(clk), .QN(n27755) );
  DFF_X2 avector10_reg_7__3_ ( .D(n24583), .CK(clk), .QN(n27754) );
  DFF_X2 avector10_reg_7__2_ ( .D(n24582), .CK(clk), .QN(n27753) );
  DFF_X2 avector10_reg_7__1_ ( .D(n24581), .CK(clk), .QN(n27752) );
  DFF_X2 avector10_reg_7__0_ ( .D(n24580), .CK(clk), .QN(n27751) );
  DFF_X2 avector10_reg_6__15_ ( .D(n24611), .CK(clk), .QN(n26998) );
  DFF_X2 avector10_reg_6__14_ ( .D(n24610), .CK(clk), .QN(n26997) );
  DFF_X2 avector10_reg_6__13_ ( .D(n24609), .CK(clk), .QN(n26996) );
  DFF_X2 avector10_reg_6__12_ ( .D(n24608), .CK(clk), .QN(n26995) );
  DFF_X2 avector10_reg_6__11_ ( .D(n24607), .CK(clk), .QN(n26994) );
  DFF_X2 avector10_reg_6__10_ ( .D(n24606), .CK(clk), .QN(n26993) );
  DFF_X2 avector10_reg_6__9_ ( .D(n24605), .CK(clk), .QN(n26992) );
  DFF_X2 avector10_reg_6__8_ ( .D(n24604), .CK(clk), .QN(n26991) );
  DFF_X2 avector10_reg_6__7_ ( .D(n24603), .CK(clk), .QN(n26990) );
  DFF_X2 avector10_reg_6__6_ ( .D(n24602), .CK(clk), .QN(n26989) );
  DFF_X2 avector10_reg_6__5_ ( .D(n24601), .CK(clk), .QN(n26988) );
  DFF_X2 avector10_reg_6__4_ ( .D(n24600), .CK(clk), .QN(n26987) );
  DFF_X2 avector10_reg_6__3_ ( .D(n24599), .CK(clk), .QN(n26986) );
  DFF_X2 avector10_reg_6__2_ ( .D(n24598), .CK(clk), .QN(n26985) );
  DFF_X2 avector10_reg_6__1_ ( .D(n24597), .CK(clk), .QN(n26984) );
  DFF_X2 avector10_reg_6__0_ ( .D(n24596), .CK(clk), .QN(n26983) );
  DFF_X2 avector10_reg_1__15_ ( .D(n24627), .CK(clk), .Q(n17577), .QN(n27254)
         );
  DFF_X2 avector10_reg_1__14_ ( .D(n24626), .CK(clk), .Q(n17614), .QN(n27253)
         );
  DFF_X2 avector10_reg_1__13_ ( .D(n24625), .CK(clk), .Q(n17651), .QN(n27252)
         );
  DFF_X2 avector10_reg_1__12_ ( .D(n24624), .CK(clk), .Q(n17688), .QN(n27251)
         );
  DFF_X2 avector10_reg_1__11_ ( .D(n24623), .CK(clk), .Q(n17725), .QN(n27250)
         );
  DFF_X2 avector10_reg_1__10_ ( .D(n24622), .CK(clk), .Q(n17762), .QN(n27249)
         );
  DFF_X2 avector10_reg_1__9_ ( .D(n24621), .CK(clk), .Q(n17799), .QN(n27248)
         );
  DFF_X2 avector10_reg_1__8_ ( .D(n24620), .CK(clk), .Q(n17836), .QN(n27247)
         );
  DFF_X2 avector10_reg_1__7_ ( .D(n24619), .CK(clk), .Q(n17873), .QN(n27246)
         );
  DFF_X2 avector10_reg_1__6_ ( .D(n24618), .CK(clk), .Q(n17910), .QN(n27245)
         );
  DFF_X2 avector10_reg_1__5_ ( .D(n24617), .CK(clk), .Q(n17947), .QN(n27244)
         );
  DFF_X2 avector10_reg_1__4_ ( .D(n24616), .CK(clk), .Q(n17984), .QN(n27243)
         );
  DFF_X2 avector10_reg_1__3_ ( .D(n24615), .CK(clk), .Q(n18021), .QN(n27242)
         );
  DFF_X2 avector10_reg_1__2_ ( .D(n24614), .CK(clk), .Q(n18058), .QN(n27241)
         );
  DFF_X2 avector10_reg_1__1_ ( .D(n24613), .CK(clk), .Q(n18095), .QN(n27240)
         );
  DFF_X2 avector10_reg_1__0_ ( .D(n24612), .CK(clk), .Q(n18132), .QN(n27239)
         );
  DFF_X2 avector10_reg_0__15_ ( .D(n24643), .CK(clk), .Q(n17578), .QN(n27510)
         );
  DFF_X2 avector10_reg_0__14_ ( .D(n24642), .CK(clk), .Q(n17615), .QN(n27509)
         );
  DFF_X2 avector10_reg_0__13_ ( .D(n24641), .CK(clk), .Q(n17652), .QN(n27508)
         );
  DFF_X2 avector10_reg_0__12_ ( .D(n24640), .CK(clk), .Q(n17689), .QN(n27507)
         );
  DFF_X2 avector10_reg_0__11_ ( .D(n24639), .CK(clk), .Q(n17726), .QN(n27506)
         );
  DFF_X2 avector10_reg_0__10_ ( .D(n24638), .CK(clk), .Q(n17763), .QN(n27505)
         );
  DFF_X2 avector10_reg_0__9_ ( .D(n24637), .CK(clk), .Q(n17800), .QN(n27504)
         );
  DFF_X2 avector10_reg_0__8_ ( .D(n24636), .CK(clk), .Q(n17837), .QN(n27503)
         );
  DFF_X2 avector10_reg_0__7_ ( .D(n24635), .CK(clk), .Q(n17874), .QN(n27502)
         );
  DFF_X2 avector10_reg_0__6_ ( .D(n24634), .CK(clk), .Q(n17911), .QN(n27501)
         );
  DFF_X2 avector10_reg_0__5_ ( .D(n24633), .CK(clk), .Q(n17948), .QN(n27500)
         );
  DFF_X2 avector10_reg_0__4_ ( .D(n24632), .CK(clk), .Q(n17985), .QN(n27499)
         );
  DFF_X2 avector10_reg_0__3_ ( .D(n24631), .CK(clk), .Q(n18022), .QN(n27498)
         );
  DFF_X2 avector10_reg_0__2_ ( .D(n24630), .CK(clk), .Q(n18059), .QN(n27497)
         );
  DFF_X2 avector10_reg_0__1_ ( .D(n24629), .CK(clk), .Q(n18096), .QN(n27496)
         );
  DFF_X2 avector10_reg_0__0_ ( .D(n24628), .CK(clk), .Q(n18133), .QN(n27495)
         );
  DFF_X2 avector03_reg_7__15_ ( .D(n23715), .CK(clk), .QN(n27590) );
  DFF_X2 avector03_reg_7__14_ ( .D(n23714), .CK(clk), .QN(n27589) );
  DFF_X2 avector03_reg_7__13_ ( .D(n23713), .CK(clk), .QN(n27588) );
  DFF_X2 avector03_reg_7__12_ ( .D(n23712), .CK(clk), .QN(n27587) );
  DFF_X2 avector03_reg_7__11_ ( .D(n23711), .CK(clk), .QN(n27586) );
  DFF_X2 avector03_reg_7__10_ ( .D(n23710), .CK(clk), .QN(n27585) );
  DFF_X2 avector03_reg_7__9_ ( .D(n23709), .CK(clk), .QN(n27584) );
  DFF_X2 avector03_reg_7__8_ ( .D(n23708), .CK(clk), .QN(n27583) );
  DFF_X2 avector03_reg_7__7_ ( .D(n23707), .CK(clk), .QN(n27582) );
  DFF_X2 avector03_reg_7__6_ ( .D(n23706), .CK(clk), .QN(n27581) );
  DFF_X2 avector03_reg_7__5_ ( .D(n23705), .CK(clk), .QN(n27580) );
  DFF_X2 avector03_reg_7__4_ ( .D(n23704), .CK(clk), .QN(n27579) );
  DFF_X2 avector03_reg_7__3_ ( .D(n23703), .CK(clk), .QN(n27578) );
  DFF_X2 avector03_reg_7__2_ ( .D(n23702), .CK(clk), .QN(n27577) );
  DFF_X2 avector03_reg_7__1_ ( .D(n23701), .CK(clk), .QN(n27576) );
  DFF_X2 avector03_reg_7__0_ ( .D(n23700), .CK(clk), .QN(n27575) );
  DFF_X2 avector03_reg_6__15_ ( .D(n23731), .CK(clk), .QN(n26822) );
  DFF_X2 avector03_reg_6__14_ ( .D(n23730), .CK(clk), .QN(n26821) );
  DFF_X2 avector03_reg_6__13_ ( .D(n23729), .CK(clk), .QN(n26820) );
  DFF_X2 avector03_reg_6__12_ ( .D(n23728), .CK(clk), .QN(n26819) );
  DFF_X2 avector03_reg_6__11_ ( .D(n23727), .CK(clk), .QN(n26818) );
  DFF_X2 avector03_reg_6__10_ ( .D(n23726), .CK(clk), .QN(n26817) );
  DFF_X2 avector03_reg_6__9_ ( .D(n23725), .CK(clk), .QN(n26816) );
  DFF_X2 avector03_reg_6__8_ ( .D(n23724), .CK(clk), .QN(n26815) );
  DFF_X2 avector03_reg_6__7_ ( .D(n23723), .CK(clk), .QN(n26814) );
  DFF_X2 avector03_reg_6__6_ ( .D(n23722), .CK(clk), .QN(n26813) );
  DFF_X2 avector03_reg_6__5_ ( .D(n23721), .CK(clk), .QN(n26812) );
  DFF_X2 avector03_reg_6__4_ ( .D(n23720), .CK(clk), .QN(n26811) );
  DFF_X2 avector03_reg_6__3_ ( .D(n23719), .CK(clk), .QN(n26810) );
  DFF_X2 avector03_reg_6__2_ ( .D(n23718), .CK(clk), .QN(n26809) );
  DFF_X2 avector03_reg_6__1_ ( .D(n23717), .CK(clk), .QN(n26808) );
  DFF_X2 avector03_reg_6__0_ ( .D(n23716), .CK(clk), .QN(n26807) );
  DFF_X2 avector03_reg_1__15_ ( .D(n23747), .CK(clk), .Q(n18178), .QN(n27078)
         );
  DFF_X2 avector03_reg_1__14_ ( .D(n23746), .CK(clk), .Q(n18215), .QN(n27077)
         );
  DFF_X2 avector03_reg_1__13_ ( .D(n23745), .CK(clk), .Q(n18252), .QN(n27076)
         );
  DFF_X2 avector03_reg_1__12_ ( .D(n23744), .CK(clk), .Q(n18289), .QN(n27075)
         );
  DFF_X2 avector03_reg_1__11_ ( .D(n23743), .CK(clk), .Q(n18326), .QN(n27074)
         );
  DFF_X2 avector03_reg_1__10_ ( .D(n23742), .CK(clk), .Q(n18363), .QN(n27073)
         );
  DFF_X2 avector03_reg_1__9_ ( .D(n23741), .CK(clk), .Q(n18400), .QN(n27072)
         );
  DFF_X2 avector03_reg_1__8_ ( .D(n23740), .CK(clk), .Q(n18437), .QN(n27071)
         );
  DFF_X2 avector03_reg_1__7_ ( .D(n23739), .CK(clk), .Q(n18474), .QN(n27070)
         );
  DFF_X2 avector03_reg_1__6_ ( .D(n23738), .CK(clk), .Q(n18511), .QN(n27069)
         );
  DFF_X2 avector03_reg_1__5_ ( .D(n23737), .CK(clk), .Q(n18548), .QN(n27068)
         );
  DFF_X2 avector03_reg_1__4_ ( .D(n23736), .CK(clk), .Q(n18585), .QN(n27067)
         );
  DFF_X2 avector03_reg_1__3_ ( .D(n23735), .CK(clk), .Q(n18622), .QN(n27066)
         );
  DFF_X2 avector03_reg_1__2_ ( .D(n23734), .CK(clk), .Q(n18659), .QN(n27065)
         );
  DFF_X2 avector03_reg_1__1_ ( .D(n23733), .CK(clk), .Q(n18696), .QN(n27064)
         );
  DFF_X2 avector03_reg_1__0_ ( .D(n23732), .CK(clk), .Q(n18733), .QN(n27063)
         );
  DFF_X2 avector03_reg_0__15_ ( .D(n23763), .CK(clk), .Q(n18179), .QN(n27334)
         );
  DFF_X2 avector03_reg_0__14_ ( .D(n23762), .CK(clk), .Q(n18216), .QN(n27333)
         );
  DFF_X2 avector03_reg_0__13_ ( .D(n23761), .CK(clk), .Q(n18253), .QN(n27332)
         );
  DFF_X2 avector03_reg_0__12_ ( .D(n23760), .CK(clk), .Q(n18290), .QN(n27331)
         );
  DFF_X2 avector03_reg_0__11_ ( .D(n23759), .CK(clk), .Q(n18327), .QN(n27330)
         );
  DFF_X2 avector03_reg_0__10_ ( .D(n23758), .CK(clk), .Q(n18364), .QN(n27329)
         );
  DFF_X2 avector03_reg_0__9_ ( .D(n23757), .CK(clk), .Q(n18401), .QN(n27328)
         );
  DFF_X2 avector03_reg_0__8_ ( .D(n23756), .CK(clk), .Q(n18438), .QN(n27327)
         );
  DFF_X2 avector03_reg_0__7_ ( .D(n23755), .CK(clk), .Q(n18475), .QN(n27326)
         );
  DFF_X2 avector03_reg_0__6_ ( .D(n23754), .CK(clk), .Q(n18512), .QN(n27325)
         );
  DFF_X2 avector03_reg_0__5_ ( .D(n23753), .CK(clk), .Q(n18549), .QN(n27324)
         );
  DFF_X2 avector03_reg_0__4_ ( .D(n23752), .CK(clk), .Q(n18586), .QN(n27323)
         );
  DFF_X2 avector03_reg_0__3_ ( .D(n23751), .CK(clk), .Q(n18623), .QN(n27322)
         );
  DFF_X2 avector03_reg_0__2_ ( .D(n23750), .CK(clk), .Q(n18660), .QN(n27321)
         );
  DFF_X2 avector03_reg_0__1_ ( .D(n23749), .CK(clk), .Q(n18697), .QN(n27320)
         );
  DFF_X2 avector03_reg_0__0_ ( .D(n23748), .CK(clk), .Q(n18734), .QN(n27319)
         );
  DFF_X2 avector02_reg_7__15_ ( .D(n24035), .CK(clk), .Q(n18157), .QN(n27654)
         );
  DFF_X2 avector02_reg_7__14_ ( .D(n24034), .CK(clk), .Q(n18194), .QN(n27653)
         );
  DFF_X2 avector02_reg_7__13_ ( .D(n24033), .CK(clk), .Q(n18231), .QN(n27652)
         );
  DFF_X2 avector02_reg_7__12_ ( .D(n24032), .CK(clk), .Q(n18268), .QN(n27651)
         );
  DFF_X2 avector02_reg_7__11_ ( .D(n24031), .CK(clk), .Q(n18305), .QN(n27650)
         );
  DFF_X2 avector02_reg_7__10_ ( .D(n24030), .CK(clk), .Q(n18342), .QN(n27649)
         );
  DFF_X2 avector02_reg_7__9_ ( .D(n24029), .CK(clk), .Q(n18379), .QN(n27648)
         );
  DFF_X2 avector02_reg_7__8_ ( .D(n24028), .CK(clk), .Q(n18416), .QN(n27647)
         );
  DFF_X2 avector02_reg_7__7_ ( .D(n24027), .CK(clk), .Q(n18453), .QN(n27646)
         );
  DFF_X2 avector02_reg_7__6_ ( .D(n24026), .CK(clk), .Q(n18490), .QN(n27645)
         );
  DFF_X2 avector02_reg_7__5_ ( .D(n24025), .CK(clk), .Q(n18527), .QN(n27644)
         );
  DFF_X2 avector02_reg_7__4_ ( .D(n24024), .CK(clk), .Q(n18564), .QN(n27643)
         );
  DFF_X2 avector02_reg_7__3_ ( .D(n24023), .CK(clk), .Q(n18601), .QN(n27642)
         );
  DFF_X2 avector02_reg_7__2_ ( .D(n24022), .CK(clk), .Q(n18638), .QN(n27641)
         );
  DFF_X2 avector02_reg_7__1_ ( .D(n24021), .CK(clk), .Q(n18675), .QN(n27640)
         );
  DFF_X2 avector02_reg_7__0_ ( .D(n24020), .CK(clk), .Q(n18712), .QN(n27639)
         );
  DFF_X2 avector02_reg_6__15_ ( .D(n24051), .CK(clk), .Q(n18155), .QN(n26886)
         );
  DFF_X2 avector02_reg_6__14_ ( .D(n24050), .CK(clk), .Q(n18192), .QN(n26885)
         );
  DFF_X2 avector02_reg_6__13_ ( .D(n24049), .CK(clk), .Q(n18229), .QN(n26884)
         );
  DFF_X2 avector02_reg_6__12_ ( .D(n24048), .CK(clk), .Q(n18266), .QN(n26883)
         );
  DFF_X2 avector02_reg_6__11_ ( .D(n24047), .CK(clk), .Q(n18303), .QN(n26882)
         );
  DFF_X2 avector02_reg_6__10_ ( .D(n24046), .CK(clk), .Q(n18340), .QN(n26881)
         );
  DFF_X2 avector02_reg_6__9_ ( .D(n24045), .CK(clk), .Q(n18377), .QN(n26880)
         );
  DFF_X2 avector02_reg_6__8_ ( .D(n24044), .CK(clk), .Q(n18414), .QN(n26879)
         );
  DFF_X2 avector02_reg_6__7_ ( .D(n24043), .CK(clk), .Q(n18451), .QN(n26878)
         );
  DFF_X2 avector02_reg_6__6_ ( .D(n24042), .CK(clk), .Q(n18488), .QN(n26877)
         );
  DFF_X2 avector02_reg_6__5_ ( .D(n24041), .CK(clk), .Q(n18525), .QN(n26876)
         );
  DFF_X2 avector02_reg_6__4_ ( .D(n24040), .CK(clk), .Q(n18562), .QN(n26875)
         );
  DFF_X2 avector02_reg_6__3_ ( .D(n24039), .CK(clk), .Q(n18599), .QN(n26874)
         );
  DFF_X2 avector02_reg_6__2_ ( .D(n24038), .CK(clk), .Q(n18636), .QN(n26873)
         );
  DFF_X2 avector02_reg_6__1_ ( .D(n24037), .CK(clk), .Q(n18673), .QN(n26872)
         );
  DFF_X2 avector02_reg_6__0_ ( .D(n24036), .CK(clk), .Q(n18710), .QN(n26871)
         );
  DFF_X2 avector02_reg_1__15_ ( .D(n24067), .CK(clk), .QN(n27142) );
  DFF_X2 avector02_reg_1__14_ ( .D(n24066), .CK(clk), .QN(n27141) );
  DFF_X2 avector02_reg_1__13_ ( .D(n24065), .CK(clk), .QN(n27140) );
  DFF_X2 avector02_reg_1__12_ ( .D(n24064), .CK(clk), .QN(n27139) );
  DFF_X2 avector02_reg_1__11_ ( .D(n24063), .CK(clk), .QN(n27138) );
  DFF_X2 avector02_reg_1__10_ ( .D(n24062), .CK(clk), .QN(n27137) );
  DFF_X2 avector02_reg_1__9_ ( .D(n24061), .CK(clk), .QN(n27136) );
  DFF_X2 avector02_reg_1__8_ ( .D(n24060), .CK(clk), .QN(n27135) );
  DFF_X2 avector02_reg_1__7_ ( .D(n24059), .CK(clk), .QN(n27134) );
  DFF_X2 avector02_reg_1__6_ ( .D(n24058), .CK(clk), .QN(n27133) );
  DFF_X2 avector02_reg_1__5_ ( .D(n24057), .CK(clk), .QN(n27132) );
  DFF_X2 avector02_reg_1__4_ ( .D(n24056), .CK(clk), .QN(n27131) );
  DFF_X2 avector02_reg_1__3_ ( .D(n24055), .CK(clk), .QN(n27130) );
  DFF_X2 avector02_reg_1__2_ ( .D(n24054), .CK(clk), .QN(n27129) );
  DFF_X2 avector02_reg_1__1_ ( .D(n24053), .CK(clk), .QN(n27128) );
  DFF_X2 avector02_reg_1__0_ ( .D(n24052), .CK(clk), .QN(n27127) );
  DFF_X2 avector02_reg_0__15_ ( .D(n24083), .CK(clk), .QN(n27398) );
  DFF_X2 avector02_reg_0__14_ ( .D(n24082), .CK(clk), .QN(n27397) );
  DFF_X2 avector02_reg_0__13_ ( .D(n24081), .CK(clk), .QN(n27396) );
  DFF_X2 avector02_reg_0__12_ ( .D(n24080), .CK(clk), .QN(n27395) );
  DFF_X2 avector02_reg_0__11_ ( .D(n24079), .CK(clk), .QN(n27394) );
  DFF_X2 avector02_reg_0__10_ ( .D(n24078), .CK(clk), .QN(n27393) );
  DFF_X2 avector02_reg_0__9_ ( .D(n24077), .CK(clk), .QN(n27392) );
  DFF_X2 avector02_reg_0__8_ ( .D(n24076), .CK(clk), .QN(n27391) );
  DFF_X2 avector02_reg_0__7_ ( .D(n24075), .CK(clk), .QN(n27390) );
  DFF_X2 avector02_reg_0__6_ ( .D(n24074), .CK(clk), .QN(n27389) );
  DFF_X2 avector02_reg_0__5_ ( .D(n24073), .CK(clk), .QN(n27388) );
  DFF_X2 avector02_reg_0__4_ ( .D(n24072), .CK(clk), .QN(n27387) );
  DFF_X2 avector02_reg_0__3_ ( .D(n24071), .CK(clk), .QN(n27386) );
  DFF_X2 avector02_reg_0__2_ ( .D(n24070), .CK(clk), .QN(n27385) );
  DFF_X2 avector02_reg_0__1_ ( .D(n24069), .CK(clk), .QN(n27384) );
  DFF_X2 avector02_reg_0__0_ ( .D(n24068), .CK(clk), .QN(n27383) );
  DFF_X2 avector01_reg_7__15_ ( .D(n24355), .CK(clk), .Q(n18166), .QN(n27718)
         );
  DFF_X2 avector01_reg_7__14_ ( .D(n24354), .CK(clk), .Q(n18203), .QN(n27717)
         );
  DFF_X2 avector01_reg_7__13_ ( .D(n24353), .CK(clk), .Q(n18240), .QN(n27716)
         );
  DFF_X2 avector01_reg_7__12_ ( .D(n24352), .CK(clk), .Q(n18277), .QN(n27715)
         );
  DFF_X2 avector01_reg_7__11_ ( .D(n24351), .CK(clk), .Q(n18314), .QN(n27714)
         );
  DFF_X2 avector01_reg_7__10_ ( .D(n24350), .CK(clk), .Q(n18351), .QN(n27713)
         );
  DFF_X2 avector01_reg_7__9_ ( .D(n24349), .CK(clk), .Q(n18388), .QN(n27712)
         );
  DFF_X2 avector01_reg_7__8_ ( .D(n24348), .CK(clk), .Q(n18425), .QN(n27711)
         );
  DFF_X2 avector01_reg_7__7_ ( .D(n24347), .CK(clk), .Q(n18462), .QN(n27710)
         );
  DFF_X2 avector01_reg_7__6_ ( .D(n24346), .CK(clk), .Q(n18499), .QN(n27709)
         );
  DFF_X2 avector01_reg_7__5_ ( .D(n24345), .CK(clk), .Q(n18536), .QN(n27708)
         );
  DFF_X2 avector01_reg_7__4_ ( .D(n24344), .CK(clk), .Q(n18573), .QN(n27707)
         );
  DFF_X2 avector01_reg_7__3_ ( .D(n24343), .CK(clk), .Q(n18610), .QN(n27706)
         );
  DFF_X2 avector01_reg_7__2_ ( .D(n24342), .CK(clk), .Q(n18647), .QN(n27705)
         );
  DFF_X2 avector01_reg_7__1_ ( .D(n24341), .CK(clk), .Q(n18684), .QN(n27704)
         );
  DFF_X2 avector01_reg_7__0_ ( .D(n24340), .CK(clk), .Q(n18721), .QN(n27703)
         );
  DFF_X2 avector01_reg_6__15_ ( .D(n24371), .CK(clk), .QN(n26950) );
  DFF_X2 avector01_reg_6__14_ ( .D(n24370), .CK(clk), .QN(n26949) );
  DFF_X2 avector01_reg_6__13_ ( .D(n24369), .CK(clk), .QN(n26948) );
  DFF_X2 avector01_reg_6__12_ ( .D(n24368), .CK(clk), .QN(n26947) );
  DFF_X2 avector01_reg_6__11_ ( .D(n24367), .CK(clk), .QN(n26946) );
  DFF_X2 avector01_reg_6__10_ ( .D(n24366), .CK(clk), .QN(n26945) );
  DFF_X2 avector01_reg_6__9_ ( .D(n24365), .CK(clk), .QN(n26944) );
  DFF_X2 avector01_reg_6__8_ ( .D(n24364), .CK(clk), .QN(n26943) );
  DFF_X2 avector01_reg_6__7_ ( .D(n24363), .CK(clk), .QN(n26942) );
  DFF_X2 avector01_reg_6__6_ ( .D(n24362), .CK(clk), .QN(n26941) );
  DFF_X2 avector01_reg_6__5_ ( .D(n24361), .CK(clk), .QN(n26940) );
  DFF_X2 avector01_reg_6__4_ ( .D(n24360), .CK(clk), .QN(n26939) );
  DFF_X2 avector01_reg_6__3_ ( .D(n24359), .CK(clk), .QN(n26938) );
  DFF_X2 avector01_reg_6__2_ ( .D(n24358), .CK(clk), .QN(n26937) );
  DFF_X2 avector01_reg_6__1_ ( .D(n24357), .CK(clk), .QN(n26936) );
  DFF_X2 avector01_reg_6__0_ ( .D(n24356), .CK(clk), .QN(n26935) );
  DFF_X2 avector01_reg_1__15_ ( .D(n24387), .CK(clk), .QN(n27206) );
  DFF_X2 avector01_reg_1__14_ ( .D(n24386), .CK(clk), .QN(n27205) );
  DFF_X2 avector01_reg_1__13_ ( .D(n24385), .CK(clk), .QN(n27204) );
  DFF_X2 avector01_reg_1__12_ ( .D(n24384), .CK(clk), .QN(n27203) );
  DFF_X2 avector01_reg_1__11_ ( .D(n24383), .CK(clk), .QN(n27202) );
  DFF_X2 avector01_reg_1__10_ ( .D(n24382), .CK(clk), .QN(n27201) );
  DFF_X2 avector01_reg_1__9_ ( .D(n24381), .CK(clk), .QN(n27200) );
  DFF_X2 avector01_reg_1__8_ ( .D(n24380), .CK(clk), .QN(n27199) );
  DFF_X2 avector01_reg_1__7_ ( .D(n24379), .CK(clk), .QN(n27198) );
  DFF_X2 avector01_reg_1__6_ ( .D(n24378), .CK(clk), .QN(n27197) );
  DFF_X2 avector01_reg_1__5_ ( .D(n24377), .CK(clk), .QN(n27196) );
  DFF_X2 avector01_reg_1__4_ ( .D(n24376), .CK(clk), .QN(n27195) );
  DFF_X2 avector01_reg_1__3_ ( .D(n24375), .CK(clk), .QN(n27194) );
  DFF_X2 avector01_reg_1__2_ ( .D(n24374), .CK(clk), .QN(n27193) );
  DFF_X2 avector01_reg_1__1_ ( .D(n24373), .CK(clk), .QN(n27192) );
  DFF_X2 avector01_reg_1__0_ ( .D(n24372), .CK(clk), .QN(n27191) );
  DFF_X2 avector01_reg_0__15_ ( .D(n24403), .CK(clk), .QN(n27462) );
  DFF_X2 avector01_reg_0__14_ ( .D(n24402), .CK(clk), .QN(n27461) );
  DFF_X2 avector01_reg_0__13_ ( .D(n24401), .CK(clk), .QN(n27460) );
  DFF_X2 avector01_reg_0__12_ ( .D(n24400), .CK(clk), .QN(n27459) );
  DFF_X2 avector01_reg_0__11_ ( .D(n24399), .CK(clk), .QN(n27458) );
  DFF_X2 avector01_reg_0__10_ ( .D(n24398), .CK(clk), .QN(n27457) );
  DFF_X2 avector01_reg_0__9_ ( .D(n24397), .CK(clk), .QN(n27456) );
  DFF_X2 avector01_reg_0__8_ ( .D(n24396), .CK(clk), .QN(n27455) );
  DFF_X2 avector01_reg_0__7_ ( .D(n24395), .CK(clk), .QN(n27454) );
  DFF_X2 avector01_reg_0__6_ ( .D(n24394), .CK(clk), .QN(n27453) );
  DFF_X2 avector01_reg_0__5_ ( .D(n24393), .CK(clk), .QN(n27452) );
  DFF_X2 avector01_reg_0__4_ ( .D(n24392), .CK(clk), .QN(n27451) );
  DFF_X2 avector01_reg_0__3_ ( .D(n24391), .CK(clk), .QN(n27450) );
  DFF_X2 avector01_reg_0__2_ ( .D(n24390), .CK(clk), .QN(n27449) );
  DFF_X2 avector01_reg_0__1_ ( .D(n24389), .CK(clk), .QN(n27448) );
  DFF_X2 avector01_reg_0__0_ ( .D(n24388), .CK(clk), .QN(n27447) );
  DFF_X2 avector00_reg_7__15_ ( .D(n24681), .CK(clk), .QN(n27782) );
  DFF_X2 avector00_reg_7__14_ ( .D(n24680), .CK(clk), .QN(n27781) );
  DFF_X2 avector00_reg_7__13_ ( .D(n24679), .CK(clk), .QN(n27780) );
  DFF_X2 avector00_reg_7__12_ ( .D(n24678), .CK(clk), .QN(n27779) );
  DFF_X2 avector00_reg_7__11_ ( .D(n24677), .CK(clk), .QN(n27778) );
  DFF_X2 avector00_reg_7__10_ ( .D(n24676), .CK(clk), .QN(n27777) );
  DFF_X2 avector00_reg_7__9_ ( .D(n24675), .CK(clk), .QN(n27776) );
  DFF_X2 avector00_reg_7__8_ ( .D(n24674), .CK(clk), .QN(n27775) );
  DFF_X2 avector00_reg_7__7_ ( .D(n24673), .CK(clk), .QN(n27774) );
  DFF_X2 avector00_reg_7__6_ ( .D(n24672), .CK(clk), .QN(n27773) );
  DFF_X2 avector00_reg_7__5_ ( .D(n24671), .CK(clk), .QN(n27772) );
  DFF_X2 avector00_reg_7__4_ ( .D(n24670), .CK(clk), .QN(n27771) );
  DFF_X2 avector00_reg_7__3_ ( .D(n24669), .CK(clk), .QN(n27770) );
  DFF_X2 avector00_reg_7__2_ ( .D(n24668), .CK(clk), .QN(n27769) );
  DFF_X2 avector00_reg_7__1_ ( .D(n24667), .CK(clk), .QN(n27768) );
  DFF_X2 avector00_reg_7__0_ ( .D(n24666), .CK(clk), .QN(n27767) );
  DFF_X2 avector00_reg_6__15_ ( .D(n24697), .CK(clk), .QN(n27014) );
  DFF_X2 avector00_reg_6__14_ ( .D(n24696), .CK(clk), .QN(n27013) );
  DFF_X2 avector00_reg_6__13_ ( .D(n24695), .CK(clk), .QN(n27012) );
  DFF_X2 avector00_reg_6__12_ ( .D(n24694), .CK(clk), .QN(n27011) );
  DFF_X2 avector00_reg_6__11_ ( .D(n24693), .CK(clk), .QN(n27010) );
  DFF_X2 avector00_reg_6__10_ ( .D(n24692), .CK(clk), .QN(n27009) );
  DFF_X2 avector00_reg_6__9_ ( .D(n24691), .CK(clk), .QN(n27008) );
  DFF_X2 avector00_reg_6__8_ ( .D(n24690), .CK(clk), .QN(n27007) );
  DFF_X2 avector00_reg_6__7_ ( .D(n24689), .CK(clk), .QN(n27006) );
  DFF_X2 avector00_reg_6__6_ ( .D(n24688), .CK(clk), .QN(n27005) );
  DFF_X2 avector00_reg_6__5_ ( .D(n24687), .CK(clk), .QN(n27004) );
  DFF_X2 avector00_reg_6__4_ ( .D(n24686), .CK(clk), .QN(n27003) );
  DFF_X2 avector00_reg_6__3_ ( .D(n24685), .CK(clk), .QN(n27002) );
  DFF_X2 avector00_reg_6__2_ ( .D(n24684), .CK(clk), .QN(n27001) );
  DFF_X2 avector00_reg_6__1_ ( .D(n24683), .CK(clk), .QN(n27000) );
  DFF_X2 avector00_reg_6__0_ ( .D(n24682), .CK(clk), .QN(n26999) );
  DFF_X2 avector00_reg_1__15_ ( .D(n24713), .CK(clk), .Q(n18169), .QN(n27270)
         );
  DFF_X2 avector00_reg_1__14_ ( .D(n24712), .CK(clk), .Q(n18206), .QN(n27269)
         );
  DFF_X2 avector00_reg_1__13_ ( .D(n24711), .CK(clk), .Q(n18243), .QN(n27268)
         );
  DFF_X2 avector00_reg_1__12_ ( .D(n24710), .CK(clk), .Q(n18280), .QN(n27267)
         );
  DFF_X2 avector00_reg_1__11_ ( .D(n24709), .CK(clk), .Q(n18317), .QN(n27266)
         );
  DFF_X2 avector00_reg_1__10_ ( .D(n24708), .CK(clk), .Q(n18354), .QN(n27265)
         );
  DFF_X2 avector00_reg_1__9_ ( .D(n24707), .CK(clk), .Q(n18391), .QN(n27264)
         );
  DFF_X2 avector00_reg_1__8_ ( .D(n24706), .CK(clk), .Q(n18428), .QN(n27263)
         );
  DFF_X2 avector00_reg_1__7_ ( .D(n24705), .CK(clk), .Q(n18465), .QN(n27262)
         );
  DFF_X2 avector00_reg_1__6_ ( .D(n24704), .CK(clk), .Q(n18502), .QN(n27261)
         );
  DFF_X2 avector00_reg_1__5_ ( .D(n24703), .CK(clk), .Q(n18539), .QN(n27260)
         );
  DFF_X2 avector00_reg_1__4_ ( .D(n24702), .CK(clk), .Q(n18576), .QN(n27259)
         );
  DFF_X2 avector00_reg_1__3_ ( .D(n24701), .CK(clk), .Q(n18613), .QN(n27258)
         );
  DFF_X2 avector00_reg_1__2_ ( .D(n24700), .CK(clk), .Q(n18650), .QN(n27257)
         );
  DFF_X2 avector00_reg_1__1_ ( .D(n24699), .CK(clk), .Q(n18687), .QN(n27256)
         );
  DFF_X2 avector00_reg_1__0_ ( .D(n24698), .CK(clk), .Q(n18724), .QN(n27255)
         );
  DFF_X2 avector00_reg_0__15_ ( .D(n24729), .CK(clk), .Q(n18170), .QN(n27526)
         );
  DFF_X2 avector00_reg_0__14_ ( .D(n24728), .CK(clk), .Q(n18207), .QN(n27525)
         );
  DFF_X2 avector00_reg_0__13_ ( .D(n24727), .CK(clk), .Q(n18244), .QN(n27524)
         );
  DFF_X2 avector00_reg_0__12_ ( .D(n24726), .CK(clk), .Q(n18281), .QN(n27523)
         );
  DFF_X2 avector00_reg_0__11_ ( .D(n24725), .CK(clk), .Q(n18318), .QN(n27522)
         );
  DFF_X2 avector00_reg_0__10_ ( .D(n24724), .CK(clk), .Q(n18355), .QN(n27521)
         );
  DFF_X2 avector00_reg_0__9_ ( .D(n24723), .CK(clk), .Q(n18392), .QN(n27520)
         );
  DFF_X2 avector00_reg_0__8_ ( .D(n24722), .CK(clk), .Q(n18429), .QN(n27519)
         );
  DFF_X2 avector00_reg_0__7_ ( .D(n24721), .CK(clk), .Q(n18466), .QN(n27518)
         );
  DFF_X2 avector00_reg_0__6_ ( .D(n24720), .CK(clk), .Q(n18503), .QN(n27517)
         );
  DFF_X2 avector00_reg_0__5_ ( .D(n24719), .CK(clk), .Q(n18540), .QN(n27516)
         );
  DFF_X2 avector00_reg_0__4_ ( .D(n24718), .CK(clk), .Q(n18577), .QN(n27515)
         );
  DFF_X2 avector00_reg_0__3_ ( .D(n24717), .CK(clk), .Q(n18614), .QN(n27514)
         );
  DFF_X2 avector00_reg_0__2_ ( .D(n24716), .CK(clk), .Q(n18651), .QN(n27513)
         );
  DFF_X2 avector00_reg_0__1_ ( .D(n24715), .CK(clk), .Q(n18688), .QN(n27512)
         );
  DFF_X2 avector00_reg_0__0_ ( .D(n24714), .CK(clk), .Q(n18725), .QN(n27511)
         );
  DFF_X2 avector33_reg_8__15_ ( .D(n23779), .CK(clk), .Q(n16407), .QN(n26582)
         );
  DFF_X2 avector33_reg_8__14_ ( .D(n23778), .CK(clk), .Q(n16444), .QN(n26581)
         );
  DFF_X2 avector33_reg_8__13_ ( .D(n23777), .CK(clk), .Q(n16481), .QN(n26580)
         );
  DFF_X2 avector33_reg_8__12_ ( .D(n23776), .CK(clk), .Q(n16518), .QN(n26579)
         );
  DFF_X2 avector33_reg_8__11_ ( .D(n23775), .CK(clk), .Q(n16555), .QN(n26578)
         );
  DFF_X2 avector33_reg_8__10_ ( .D(n23774), .CK(clk), .Q(n16592), .QN(n26577)
         );
  DFF_X2 avector33_reg_8__9_ ( .D(n23773), .CK(clk), .Q(n16629), .QN(n26576)
         );
  DFF_X2 avector33_reg_8__8_ ( .D(n23772), .CK(clk), .Q(n16666), .QN(n26575)
         );
  DFF_X2 avector33_reg_8__7_ ( .D(n23771), .CK(clk), .Q(n16703), .QN(n26574)
         );
  DFF_X2 avector33_reg_8__6_ ( .D(n23770), .CK(clk), .Q(n16740), .QN(n26573)
         );
  DFF_X2 avector33_reg_8__5_ ( .D(n23769), .CK(clk), .Q(n16777), .QN(n26572)
         );
  DFF_X2 avector33_reg_8__4_ ( .D(n23768), .CK(clk), .Q(n16814), .QN(n26571)
         );
  DFF_X2 avector33_reg_8__3_ ( .D(n23767), .CK(clk), .Q(n16851), .QN(n26570)
         );
  DFF_X2 avector33_reg_8__2_ ( .D(n23766), .CK(clk), .Q(n16888), .QN(n26569)
         );
  DFF_X2 avector33_reg_8__1_ ( .D(n23765), .CK(clk), .Q(n16925), .QN(n26568)
         );
  DFF_X2 avector33_reg_8__0_ ( .D(n23764), .CK(clk), .Q(n16962), .QN(n26567)
         );
  DFF_X2 bvector3_reg_8__3_ ( .D(n23354), .CK(clk), .Q(n18899), .QN(n27817) );
  DFF_X2 bvector3_reg_8__2_ ( .D(n23353), .CK(clk), .Q(n18862), .QN(n27816) );
  DFF_X2 bvector3_reg_8__0_ ( .D(n23351), .CK(clk), .Q(n18788), .QN(n27814) );
  DFF_X2 bvector2_reg_8__3_ ( .D(n23107), .CK(clk), .QN(n28057) );
  DFF_X2 bvector2_reg_8__2_ ( .D(n23106), .CK(clk), .QN(n28056) );
  DFF_X2 bvector2_reg_8__0_ ( .D(n23104), .CK(clk), .QN(n28054) );
  DFF_X2 bvector1_reg_8__3_ ( .D(n23187), .CK(clk), .Q(n18881), .QN(n27977) );
  DFF_X2 bvector1_reg_8__2_ ( .D(n23186), .CK(clk), .Q(n18844), .QN(n27976) );
  DFF_X2 bvector1_reg_8__0_ ( .D(n23184), .CK(clk), .Q(n18770), .QN(n27974) );
  DFF_X2 bvector0_reg_8__3_ ( .D(n23274), .CK(clk), .QN(n27897) );
  DFF_X2 bvector0_reg_8__2_ ( .D(n23273), .CK(clk), .QN(n27896) );
  DFF_X2 bvector0_reg_8__0_ ( .D(n23271), .CK(clk), .QN(n27894) );
  DFF_X2 bvector3_reg_7__3_ ( .D(n23370), .CK(clk), .QN(n27833) );
  DFF_X2 bvector3_reg_7__2_ ( .D(n23369), .CK(clk), .QN(n27832) );
  DFF_X2 bvector3_reg_7__0_ ( .D(n23367), .CK(clk), .QN(n27830) );
  DFF_X2 bvector3_reg_6__3_ ( .D(n23386), .CK(clk), .Q(n18898), .QN(n27849) );
  DFF_X2 bvector3_reg_6__2_ ( .D(n23385), .CK(clk), .Q(n18861), .QN(n27848) );
  DFF_X2 bvector3_reg_6__0_ ( .D(n23383), .CK(clk), .Q(n18787), .QN(n27846) );
  DFF_X2 bvector3_reg_1__3_ ( .D(n23402), .CK(clk), .QN(n27865) );
  DFF_X2 bvector3_reg_1__2_ ( .D(n23401), .CK(clk), .QN(n27864) );
  DFF_X2 bvector3_reg_1__0_ ( .D(n23399), .CK(clk), .QN(n27862) );
  DFF_X2 bvector3_reg_0__3_ ( .D(n23418), .CK(clk), .QN(n27881) );
  DFF_X2 bvector3_reg_0__2_ ( .D(n23417), .CK(clk), .QN(n27880) );
  DFF_X2 bvector3_reg_0__0_ ( .D(n23415), .CK(clk), .QN(n27878) );
  DFF_X2 bvector2_reg_7__3_ ( .D(n23123), .CK(clk), .QN(n28073) );
  DFF_X2 bvector2_reg_7__2_ ( .D(n23122), .CK(clk), .QN(n28072) );
  DFF_X2 bvector2_reg_7__0_ ( .D(n23120), .CK(clk), .QN(n28070) );
  DFF_X2 bvector2_reg_6__3_ ( .D(n23139), .CK(clk), .QN(n28089) );
  DFF_X2 bvector2_reg_6__2_ ( .D(n23138), .CK(clk), .QN(n28088) );
  DFF_X2 bvector2_reg_6__0_ ( .D(n23136), .CK(clk), .QN(n28086) );
  DFF_X2 bvector2_reg_1__3_ ( .D(n23155), .CK(clk), .Q(n18867), .QN(n28105) );
  DFF_X2 bvector2_reg_1__2_ ( .D(n23154), .CK(clk), .Q(n18830), .QN(n28104) );
  DFF_X2 bvector2_reg_1__0_ ( .D(n23152), .CK(clk), .Q(n18756), .QN(n28102) );
  DFF_X2 bvector2_reg_0__3_ ( .D(n23171), .CK(clk), .Q(n18868), .QN(n28121) );
  DFF_X2 bvector2_reg_0__2_ ( .D(n23170), .CK(clk), .Q(n18831), .QN(n28120) );
  DFF_X2 bvector2_reg_0__0_ ( .D(n23168), .CK(clk), .Q(n18757), .QN(n28118) );
  DFF_X2 bvector1_reg_7__3_ ( .D(n23203), .CK(clk), .Q(n18882), .QN(n27993) );
  DFF_X2 bvector1_reg_7__2_ ( .D(n23202), .CK(clk), .Q(n18845), .QN(n27992) );
  DFF_X2 bvector1_reg_7__0_ ( .D(n23200), .CK(clk), .Q(n18771), .QN(n27990) );
  DFF_X2 bvector1_reg_6__3_ ( .D(n23219), .CK(clk), .QN(n28009) );
  DFF_X2 bvector1_reg_6__2_ ( .D(n23218), .CK(clk), .QN(n28008) );
  DFF_X2 bvector1_reg_6__0_ ( .D(n23216), .CK(clk), .QN(n28006) );
  DFF_X2 bvector1_reg_1__3_ ( .D(n23235), .CK(clk), .Q(n18876), .QN(n28025) );
  DFF_X2 bvector1_reg_1__2_ ( .D(n23234), .CK(clk), .Q(n18839), .QN(n28024) );
  DFF_X2 bvector1_reg_1__0_ ( .D(n23232), .CK(clk), .Q(n18765), .QN(n28022) );
  DFF_X2 bvector1_reg_0__3_ ( .D(n23251), .CK(clk), .Q(n18877), .QN(n28041) );
  DFF_X2 bvector1_reg_0__2_ ( .D(n23250), .CK(clk), .Q(n18840), .QN(n28040) );
  DFF_X2 bvector1_reg_0__0_ ( .D(n23248), .CK(clk), .Q(n18766), .QN(n28038) );
  DFF_X2 bvector0_reg_7__3_ ( .D(n23290), .CK(clk), .QN(n27913) );
  DFF_X2 bvector0_reg_7__2_ ( .D(n23289), .CK(clk), .QN(n27912) );
  DFF_X2 bvector0_reg_7__0_ ( .D(n23287), .CK(clk), .QN(n27910) );
  DFF_X2 bvector0_reg_6__3_ ( .D(n23306), .CK(clk), .QN(n27929) );
  DFF_X2 bvector0_reg_6__2_ ( .D(n23305), .CK(clk), .QN(n27928) );
  DFF_X2 bvector0_reg_6__0_ ( .D(n23303), .CK(clk), .QN(n27926) );
  DFF_X2 bvector0_reg_1__3_ ( .D(n23322), .CK(clk), .QN(n27945) );
  DFF_X2 bvector0_reg_1__2_ ( .D(n23321), .CK(clk), .QN(n27944) );
  DFF_X2 bvector0_reg_1__0_ ( .D(n23319), .CK(clk), .QN(n27942) );
  DFF_X2 bvector0_reg_0__3_ ( .D(n23338), .CK(clk), .QN(n27961) );
  DFF_X2 bvector0_reg_0__2_ ( .D(n23337), .CK(clk), .QN(n27960) );
  DFF_X2 bvector0_reg_0__0_ ( .D(n23335), .CK(clk), .QN(n27958) );
  DFF_X2 bvector3_reg_8__1_ ( .D(n23352), .CK(clk), .Q(n18825), .QN(n27815) );
  DFF_X2 bvector2_reg_8__1_ ( .D(n23105), .CK(clk), .QN(n28055) );
  DFF_X2 bvector1_reg_8__1_ ( .D(n23185), .CK(clk), .Q(n18807), .QN(n27975) );
  DFF_X2 bvector0_reg_8__1_ ( .D(n23272), .CK(clk), .QN(n27895) );
  DFF_X2 bvector3_reg_7__1_ ( .D(n23368), .CK(clk), .QN(n27831) );
  DFF_X2 bvector3_reg_6__1_ ( .D(n23384), .CK(clk), .Q(n18824), .QN(n27847) );
  DFF_X2 bvector3_reg_1__1_ ( .D(n23400), .CK(clk), .QN(n27863) );
  DFF_X2 bvector3_reg_0__1_ ( .D(n23416), .CK(clk), .QN(n27879) );
  DFF_X2 bvector2_reg_7__1_ ( .D(n23121), .CK(clk), .QN(n28071) );
  DFF_X2 bvector2_reg_6__1_ ( .D(n23137), .CK(clk), .QN(n28087) );
  DFF_X2 bvector2_reg_1__1_ ( .D(n23153), .CK(clk), .Q(n18793), .QN(n28103) );
  DFF_X2 bvector2_reg_0__1_ ( .D(n23169), .CK(clk), .Q(n18794), .QN(n28119) );
  DFF_X2 bvector1_reg_7__1_ ( .D(n23201), .CK(clk), .Q(n18808), .QN(n27991) );
  DFF_X2 bvector1_reg_6__1_ ( .D(n23217), .CK(clk), .QN(n28007) );
  DFF_X2 bvector1_reg_1__1_ ( .D(n23233), .CK(clk), .Q(n18802), .QN(n28023) );
  DFF_X2 bvector1_reg_0__1_ ( .D(n23249), .CK(clk), .Q(n18803), .QN(n28039) );
  DFF_X2 bvector0_reg_7__1_ ( .D(n23288), .CK(clk), .QN(n27911) );
  DFF_X2 bvector0_reg_6__1_ ( .D(n23304), .CK(clk), .QN(n27927) );
  DFF_X2 bvector0_reg_1__1_ ( .D(n23320), .CK(clk), .QN(n27943) );
  DFF_X2 bvector0_reg_0__1_ ( .D(n23336), .CK(clk), .QN(n27959) );
  DFF_X2 bvector3_reg_8__15_ ( .D(n23366), .CK(clk), .Q(n19343), .QN(n27829)
         );
  DFF_X2 bvector3_reg_8__14_ ( .D(n23365), .CK(clk), .Q(n19306), .QN(n27828)
         );
  DFF_X2 bvector3_reg_8__13_ ( .D(n23364), .CK(clk), .Q(n19269), .QN(n27827)
         );
  DFF_X2 bvector3_reg_8__12_ ( .D(n23363), .CK(clk), .Q(n19232), .QN(n27826)
         );
  DFF_X2 bvector3_reg_8__11_ ( .D(n23362), .CK(clk), .Q(n19195), .QN(n27825)
         );
  DFF_X2 bvector3_reg_8__10_ ( .D(n23361), .CK(clk), .Q(n19158), .QN(n27824)
         );
  DFF_X2 bvector3_reg_8__9_ ( .D(n23360), .CK(clk), .Q(n19121), .QN(n27823) );
  DFF_X2 bvector3_reg_8__8_ ( .D(n23359), .CK(clk), .Q(n19084), .QN(n27822) );
  DFF_X2 bvector3_reg_8__7_ ( .D(n23358), .CK(clk), .Q(n19047), .QN(n27821) );
  DFF_X2 bvector3_reg_8__6_ ( .D(n23357), .CK(clk), .Q(n19010), .QN(n27820) );
  DFF_X2 bvector3_reg_8__5_ ( .D(n23356), .CK(clk), .Q(n18973), .QN(n27819) );
  DFF_X2 bvector3_reg_8__4_ ( .D(n23355), .CK(clk), .Q(n18936), .QN(n27818) );
  DFF_X2 bvector2_reg_8__15_ ( .D(n23119), .CK(clk), .QN(n28069) );
  DFF_X2 bvector2_reg_8__14_ ( .D(n23118), .CK(clk), .QN(n28068) );
  DFF_X2 bvector2_reg_8__13_ ( .D(n23117), .CK(clk), .QN(n28067) );
  DFF_X2 bvector2_reg_8__12_ ( .D(n23116), .CK(clk), .QN(n28066) );
  DFF_X2 bvector2_reg_8__11_ ( .D(n23115), .CK(clk), .QN(n28065) );
  DFF_X2 bvector2_reg_8__10_ ( .D(n23114), .CK(clk), .QN(n28064) );
  DFF_X2 bvector2_reg_8__9_ ( .D(n23113), .CK(clk), .QN(n28063) );
  DFF_X2 bvector2_reg_8__8_ ( .D(n23112), .CK(clk), .QN(n28062) );
  DFF_X2 bvector2_reg_8__7_ ( .D(n23111), .CK(clk), .QN(n28061) );
  DFF_X2 bvector2_reg_8__6_ ( .D(n23110), .CK(clk), .QN(n28060) );
  DFF_X2 bvector2_reg_8__5_ ( .D(n23109), .CK(clk), .QN(n28059) );
  DFF_X2 bvector2_reg_8__4_ ( .D(n23108), .CK(clk), .QN(n28058) );
  DFF_X2 bvector1_reg_8__15_ ( .D(n23199), .CK(clk), .Q(n19325), .QN(n27989)
         );
  DFF_X2 bvector1_reg_8__14_ ( .D(n23198), .CK(clk), .Q(n19288), .QN(n27988)
         );
  DFF_X2 bvector1_reg_8__13_ ( .D(n23197), .CK(clk), .Q(n19251), .QN(n27987)
         );
  DFF_X2 bvector1_reg_8__12_ ( .D(n23196), .CK(clk), .Q(n19214), .QN(n27986)
         );
  DFF_X2 bvector1_reg_8__11_ ( .D(n23195), .CK(clk), .Q(n19177), .QN(n27985)
         );
  DFF_X2 bvector1_reg_8__10_ ( .D(n23194), .CK(clk), .Q(n19140), .QN(n27984)
         );
  DFF_X2 bvector1_reg_8__9_ ( .D(n23193), .CK(clk), .Q(n19103), .QN(n27983) );
  DFF_X2 bvector1_reg_8__8_ ( .D(n23192), .CK(clk), .Q(n19066), .QN(n27982) );
  DFF_X2 bvector1_reg_8__7_ ( .D(n23191), .CK(clk), .Q(n19029), .QN(n27981) );
  DFF_X2 bvector1_reg_8__6_ ( .D(n23190), .CK(clk), .Q(n18992), .QN(n27980) );
  DFF_X2 bvector1_reg_8__5_ ( .D(n23189), .CK(clk), .Q(n18955), .QN(n27979) );
  DFF_X2 bvector1_reg_8__4_ ( .D(n23188), .CK(clk), .Q(n18918), .QN(n27978) );
  DFF_X2 bvector0_reg_8__15_ ( .D(n23286), .CK(clk), .QN(n27909) );
  DFF_X2 bvector0_reg_8__14_ ( .D(n23285), .CK(clk), .QN(n27908) );
  DFF_X2 bvector0_reg_8__13_ ( .D(n23284), .CK(clk), .QN(n27907) );
  DFF_X2 bvector0_reg_8__12_ ( .D(n23283), .CK(clk), .QN(n27906) );
  DFF_X2 bvector0_reg_8__11_ ( .D(n23282), .CK(clk), .QN(n27905) );
  DFF_X2 bvector0_reg_8__10_ ( .D(n23281), .CK(clk), .QN(n27904) );
  DFF_X2 bvector0_reg_8__9_ ( .D(n23280), .CK(clk), .QN(n27903) );
  DFF_X2 bvector0_reg_8__8_ ( .D(n23279), .CK(clk), .QN(n27902) );
  DFF_X2 bvector0_reg_8__7_ ( .D(n23278), .CK(clk), .QN(n27901) );
  DFF_X2 bvector0_reg_8__6_ ( .D(n23277), .CK(clk), .QN(n27900) );
  DFF_X2 bvector0_reg_8__5_ ( .D(n23276), .CK(clk), .QN(n27899) );
  DFF_X2 bvector0_reg_8__4_ ( .D(n23275), .CK(clk), .QN(n27898) );
  DFF_X2 bvector3_reg_7__15_ ( .D(n23382), .CK(clk), .QN(n27845) );
  DFF_X2 bvector3_reg_7__14_ ( .D(n23381), .CK(clk), .QN(n27844) );
  DFF_X2 bvector3_reg_7__13_ ( .D(n23380), .CK(clk), .QN(n27843) );
  DFF_X2 bvector3_reg_7__12_ ( .D(n23379), .CK(clk), .QN(n27842) );
  DFF_X2 bvector3_reg_7__11_ ( .D(n23378), .CK(clk), .QN(n27841) );
  DFF_X2 bvector3_reg_7__10_ ( .D(n23377), .CK(clk), .QN(n27840) );
  DFF_X2 bvector3_reg_7__9_ ( .D(n23376), .CK(clk), .QN(n27839) );
  DFF_X2 bvector3_reg_7__8_ ( .D(n23375), .CK(clk), .QN(n27838) );
  DFF_X2 bvector3_reg_7__7_ ( .D(n23374), .CK(clk), .QN(n27837) );
  DFF_X2 bvector3_reg_7__6_ ( .D(n23373), .CK(clk), .QN(n27836) );
  DFF_X2 bvector3_reg_7__5_ ( .D(n23372), .CK(clk), .QN(n27835) );
  DFF_X2 bvector3_reg_7__4_ ( .D(n23371), .CK(clk), .QN(n27834) );
  DFF_X2 bvector3_reg_6__15_ ( .D(n23398), .CK(clk), .Q(n19342), .QN(n27861)
         );
  DFF_X2 bvector3_reg_6__14_ ( .D(n23397), .CK(clk), .Q(n19305), .QN(n27860)
         );
  DFF_X2 bvector3_reg_6__13_ ( .D(n23396), .CK(clk), .Q(n19268), .QN(n27859)
         );
  DFF_X2 bvector3_reg_6__12_ ( .D(n23395), .CK(clk), .Q(n19231), .QN(n27858)
         );
  DFF_X2 bvector3_reg_6__11_ ( .D(n23394), .CK(clk), .Q(n19194), .QN(n27857)
         );
  DFF_X2 bvector3_reg_6__10_ ( .D(n23393), .CK(clk), .Q(n19157), .QN(n27856)
         );
  DFF_X2 bvector3_reg_6__9_ ( .D(n23392), .CK(clk), .Q(n19120), .QN(n27855) );
  DFF_X2 bvector3_reg_6__8_ ( .D(n23391), .CK(clk), .Q(n19083), .QN(n27854) );
  DFF_X2 bvector3_reg_6__7_ ( .D(n23390), .CK(clk), .Q(n19046), .QN(n27853) );
  DFF_X2 bvector3_reg_6__6_ ( .D(n23389), .CK(clk), .Q(n19009), .QN(n27852) );
  DFF_X2 bvector3_reg_6__5_ ( .D(n23388), .CK(clk), .Q(n18972), .QN(n27851) );
  DFF_X2 bvector3_reg_6__4_ ( .D(n23387), .CK(clk), .Q(n18935), .QN(n27850) );
  DFF_X2 bvector3_reg_1__15_ ( .D(n23414), .CK(clk), .QN(n27877) );
  DFF_X2 bvector3_reg_1__14_ ( .D(n23413), .CK(clk), .QN(n27876) );
  DFF_X2 bvector3_reg_1__13_ ( .D(n23412), .CK(clk), .QN(n27875) );
  DFF_X2 bvector3_reg_1__12_ ( .D(n23411), .CK(clk), .QN(n27874) );
  DFF_X2 bvector3_reg_1__11_ ( .D(n23410), .CK(clk), .QN(n27873) );
  DFF_X2 bvector3_reg_1__10_ ( .D(n23409), .CK(clk), .QN(n27872) );
  DFF_X2 bvector3_reg_1__9_ ( .D(n23408), .CK(clk), .QN(n27871) );
  DFF_X2 bvector3_reg_1__8_ ( .D(n23407), .CK(clk), .QN(n27870) );
  DFF_X2 bvector3_reg_1__7_ ( .D(n23406), .CK(clk), .QN(n27869) );
  DFF_X2 bvector3_reg_1__6_ ( .D(n23405), .CK(clk), .QN(n27868) );
  DFF_X2 bvector3_reg_1__5_ ( .D(n23404), .CK(clk), .QN(n27867) );
  DFF_X2 bvector3_reg_1__4_ ( .D(n23403), .CK(clk), .QN(n27866) );
  DFF_X2 bvector3_reg_0__15_ ( .D(n23430), .CK(clk), .QN(n27893) );
  DFF_X2 bvector3_reg_0__14_ ( .D(n23429), .CK(clk), .QN(n27892) );
  DFF_X2 bvector3_reg_0__13_ ( .D(n23428), .CK(clk), .QN(n27891) );
  DFF_X2 bvector3_reg_0__12_ ( .D(n23427), .CK(clk), .QN(n27890) );
  DFF_X2 bvector3_reg_0__11_ ( .D(n23426), .CK(clk), .QN(n27889) );
  DFF_X2 bvector3_reg_0__10_ ( .D(n23425), .CK(clk), .QN(n27888) );
  DFF_X2 bvector3_reg_0__9_ ( .D(n23424), .CK(clk), .QN(n27887) );
  DFF_X2 bvector3_reg_0__8_ ( .D(n23423), .CK(clk), .QN(n27886) );
  DFF_X2 bvector3_reg_0__7_ ( .D(n23422), .CK(clk), .QN(n27885) );
  DFF_X2 bvector3_reg_0__6_ ( .D(n23421), .CK(clk), .QN(n27884) );
  DFF_X2 bvector3_reg_0__5_ ( .D(n23420), .CK(clk), .QN(n27883) );
  DFF_X2 bvector3_reg_0__4_ ( .D(n23419), .CK(clk), .QN(n27882) );
  DFF_X2 bvector2_reg_7__15_ ( .D(n23135), .CK(clk), .QN(n28085) );
  DFF_X2 bvector2_reg_7__14_ ( .D(n23134), .CK(clk), .QN(n28084) );
  DFF_X2 bvector2_reg_7__13_ ( .D(n23133), .CK(clk), .QN(n28083) );
  DFF_X2 bvector2_reg_7__12_ ( .D(n23132), .CK(clk), .QN(n28082) );
  DFF_X2 bvector2_reg_7__11_ ( .D(n23131), .CK(clk), .QN(n28081) );
  DFF_X2 bvector2_reg_7__10_ ( .D(n23130), .CK(clk), .QN(n28080) );
  DFF_X2 bvector2_reg_7__9_ ( .D(n23129), .CK(clk), .QN(n28079) );
  DFF_X2 bvector2_reg_7__8_ ( .D(n23128), .CK(clk), .QN(n28078) );
  DFF_X2 bvector2_reg_7__7_ ( .D(n23127), .CK(clk), .QN(n28077) );
  DFF_X2 bvector2_reg_7__6_ ( .D(n23126), .CK(clk), .QN(n28076) );
  DFF_X2 bvector2_reg_7__5_ ( .D(n23125), .CK(clk), .QN(n28075) );
  DFF_X2 bvector2_reg_7__4_ ( .D(n23124), .CK(clk), .QN(n28074) );
  DFF_X2 bvector2_reg_6__15_ ( .D(n23151), .CK(clk), .QN(n28101) );
  DFF_X2 bvector2_reg_6__14_ ( .D(n23150), .CK(clk), .QN(n28100) );
  DFF_X2 bvector2_reg_6__13_ ( .D(n23149), .CK(clk), .QN(n28099) );
  DFF_X2 bvector2_reg_6__12_ ( .D(n23148), .CK(clk), .QN(n28098) );
  DFF_X2 bvector2_reg_6__11_ ( .D(n23147), .CK(clk), .QN(n28097) );
  DFF_X2 bvector2_reg_6__10_ ( .D(n23146), .CK(clk), .QN(n28096) );
  DFF_X2 bvector2_reg_6__9_ ( .D(n23145), .CK(clk), .QN(n28095) );
  DFF_X2 bvector2_reg_6__8_ ( .D(n23144), .CK(clk), .QN(n28094) );
  DFF_X2 bvector2_reg_6__7_ ( .D(n23143), .CK(clk), .QN(n28093) );
  DFF_X2 bvector2_reg_6__6_ ( .D(n23142), .CK(clk), .QN(n28092) );
  DFF_X2 bvector2_reg_6__5_ ( .D(n23141), .CK(clk), .QN(n28091) );
  DFF_X2 bvector2_reg_6__4_ ( .D(n23140), .CK(clk), .QN(n28090) );
  DFF_X2 bvector2_reg_1__15_ ( .D(n23167), .CK(clk), .Q(n19311), .QN(n28117)
         );
  DFF_X2 bvector2_reg_1__14_ ( .D(n23166), .CK(clk), .Q(n19274), .QN(n28116)
         );
  DFF_X2 bvector2_reg_1__13_ ( .D(n23165), .CK(clk), .Q(n19237), .QN(n28115)
         );
  DFF_X2 bvector2_reg_1__12_ ( .D(n23164), .CK(clk), .Q(n19200), .QN(n28114)
         );
  DFF_X2 bvector2_reg_1__11_ ( .D(n23163), .CK(clk), .Q(n19163), .QN(n28113)
         );
  DFF_X2 bvector2_reg_1__10_ ( .D(n23162), .CK(clk), .Q(n19126), .QN(n28112)
         );
  DFF_X2 bvector2_reg_1__9_ ( .D(n23161), .CK(clk), .Q(n19089), .QN(n28111) );
  DFF_X2 bvector2_reg_1__8_ ( .D(n23160), .CK(clk), .Q(n19052), .QN(n28110) );
  DFF_X2 bvector2_reg_1__7_ ( .D(n23159), .CK(clk), .Q(n19015), .QN(n28109) );
  DFF_X2 bvector2_reg_1__6_ ( .D(n23158), .CK(clk), .Q(n18978), .QN(n28108) );
  DFF_X2 bvector2_reg_1__5_ ( .D(n23157), .CK(clk), .Q(n18941), .QN(n28107) );
  DFF_X2 bvector2_reg_1__4_ ( .D(n23156), .CK(clk), .Q(n18904), .QN(n28106) );
  DFF_X2 bvector2_reg_0__15_ ( .D(n23183), .CK(clk), .Q(n19312), .QN(n28133)
         );
  DFF_X2 bvector2_reg_0__14_ ( .D(n23182), .CK(clk), .Q(n19275), .QN(n28132)
         );
  DFF_X2 bvector2_reg_0__13_ ( .D(n23181), .CK(clk), .Q(n19238), .QN(n28131)
         );
  DFF_X2 bvector2_reg_0__12_ ( .D(n23180), .CK(clk), .Q(n19201), .QN(n28130)
         );
  DFF_X2 bvector2_reg_0__11_ ( .D(n23179), .CK(clk), .Q(n19164), .QN(n28129)
         );
  DFF_X2 bvector2_reg_0__10_ ( .D(n23178), .CK(clk), .Q(n19127), .QN(n28128)
         );
  DFF_X2 bvector2_reg_0__9_ ( .D(n23177), .CK(clk), .Q(n19090), .QN(n28127) );
  DFF_X2 bvector2_reg_0__8_ ( .D(n23176), .CK(clk), .Q(n19053), .QN(n28126) );
  DFF_X2 bvector2_reg_0__7_ ( .D(n23175), .CK(clk), .Q(n19016), .QN(n28125) );
  DFF_X2 bvector2_reg_0__6_ ( .D(n23174), .CK(clk), .Q(n18979), .QN(n28124) );
  DFF_X2 bvector2_reg_0__5_ ( .D(n23173), .CK(clk), .Q(n18942), .QN(n28123) );
  DFF_X2 bvector2_reg_0__4_ ( .D(n23172), .CK(clk), .Q(n18905), .QN(n28122) );
  DFF_X2 bvector1_reg_7__15_ ( .D(n23215), .CK(clk), .Q(n19326), .QN(n28005)
         );
  DFF_X2 bvector1_reg_7__14_ ( .D(n23214), .CK(clk), .Q(n19289), .QN(n28004)
         );
  DFF_X2 bvector1_reg_7__13_ ( .D(n23213), .CK(clk), .Q(n19252), .QN(n28003)
         );
  DFF_X2 bvector1_reg_7__12_ ( .D(n23212), .CK(clk), .Q(n19215), .QN(n28002)
         );
  DFF_X2 bvector1_reg_7__11_ ( .D(n23211), .CK(clk), .Q(n19178), .QN(n28001)
         );
  DFF_X2 bvector1_reg_7__10_ ( .D(n23210), .CK(clk), .Q(n19141), .QN(n28000)
         );
  DFF_X2 bvector1_reg_7__9_ ( .D(n23209), .CK(clk), .Q(n19104), .QN(n27999) );
  DFF_X2 bvector1_reg_7__8_ ( .D(n23208), .CK(clk), .Q(n19067), .QN(n27998) );
  DFF_X2 bvector1_reg_7__7_ ( .D(n23207), .CK(clk), .Q(n19030), .QN(n27997) );
  DFF_X2 bvector1_reg_7__6_ ( .D(n23206), .CK(clk), .Q(n18993), .QN(n27996) );
  DFF_X2 bvector1_reg_7__5_ ( .D(n23205), .CK(clk), .Q(n18956), .QN(n27995) );
  DFF_X2 bvector1_reg_7__4_ ( .D(n23204), .CK(clk), .Q(n18919), .QN(n27994) );
  DFF_X2 bvector1_reg_6__15_ ( .D(n23231), .CK(clk), .QN(n28021) );
  DFF_X2 bvector1_reg_6__14_ ( .D(n23230), .CK(clk), .QN(n28020) );
  DFF_X2 bvector1_reg_6__13_ ( .D(n23229), .CK(clk), .QN(n28019) );
  DFF_X2 bvector1_reg_6__12_ ( .D(n23228), .CK(clk), .QN(n28018) );
  DFF_X2 bvector1_reg_6__11_ ( .D(n23227), .CK(clk), .QN(n28017) );
  DFF_X2 bvector1_reg_6__10_ ( .D(n23226), .CK(clk), .QN(n28016) );
  DFF_X2 bvector1_reg_6__9_ ( .D(n23225), .CK(clk), .QN(n28015) );
  DFF_X2 bvector1_reg_6__8_ ( .D(n23224), .CK(clk), .QN(n28014) );
  DFF_X2 bvector1_reg_6__7_ ( .D(n23223), .CK(clk), .QN(n28013) );
  DFF_X2 bvector1_reg_6__6_ ( .D(n23222), .CK(clk), .QN(n28012) );
  DFF_X2 bvector1_reg_6__5_ ( .D(n23221), .CK(clk), .QN(n28011) );
  DFF_X2 bvector1_reg_6__4_ ( .D(n23220), .CK(clk), .QN(n28010) );
  DFF_X2 bvector1_reg_1__15_ ( .D(n23247), .CK(clk), .Q(n19320), .QN(n28037)
         );
  DFF_X2 bvector1_reg_1__14_ ( .D(n23246), .CK(clk), .Q(n19283), .QN(n28036)
         );
  DFF_X2 bvector1_reg_1__13_ ( .D(n23245), .CK(clk), .Q(n19246), .QN(n28035)
         );
  DFF_X2 bvector1_reg_1__12_ ( .D(n23244), .CK(clk), .Q(n19209), .QN(n28034)
         );
  DFF_X2 bvector1_reg_1__11_ ( .D(n23243), .CK(clk), .Q(n19172), .QN(n28033)
         );
  DFF_X2 bvector1_reg_1__10_ ( .D(n23242), .CK(clk), .Q(n19135), .QN(n28032)
         );
  DFF_X2 bvector1_reg_1__9_ ( .D(n23241), .CK(clk), .Q(n19098), .QN(n28031) );
  DFF_X2 bvector1_reg_1__8_ ( .D(n23240), .CK(clk), .Q(n19061), .QN(n28030) );
  DFF_X2 bvector1_reg_1__7_ ( .D(n23239), .CK(clk), .Q(n19024), .QN(n28029) );
  DFF_X2 bvector1_reg_1__6_ ( .D(n23238), .CK(clk), .Q(n18987), .QN(n28028) );
  DFF_X2 bvector1_reg_1__5_ ( .D(n23237), .CK(clk), .Q(n18950), .QN(n28027) );
  DFF_X2 bvector1_reg_1__4_ ( .D(n23236), .CK(clk), .Q(n18913), .QN(n28026) );
  DFF_X2 bvector1_reg_0__15_ ( .D(n23263), .CK(clk), .Q(n19321), .QN(n28053)
         );
  DFF_X2 bvector1_reg_0__14_ ( .D(n23262), .CK(clk), .Q(n19284), .QN(n28052)
         );
  DFF_X2 bvector1_reg_0__13_ ( .D(n23261), .CK(clk), .Q(n19247), .QN(n28051)
         );
  DFF_X2 bvector1_reg_0__12_ ( .D(n23260), .CK(clk), .Q(n19210), .QN(n28050)
         );
  DFF_X2 bvector1_reg_0__11_ ( .D(n23259), .CK(clk), .Q(n19173), .QN(n28049)
         );
  DFF_X2 bvector1_reg_0__10_ ( .D(n23258), .CK(clk), .Q(n19136), .QN(n28048)
         );
  DFF_X2 bvector1_reg_0__9_ ( .D(n23257), .CK(clk), .Q(n19099), .QN(n28047) );
  DFF_X2 bvector1_reg_0__8_ ( .D(n23256), .CK(clk), .Q(n19062), .QN(n28046) );
  DFF_X2 bvector1_reg_0__7_ ( .D(n23255), .CK(clk), .Q(n19025), .QN(n28045) );
  DFF_X2 bvector1_reg_0__6_ ( .D(n23254), .CK(clk), .Q(n18988), .QN(n28044) );
  DFF_X2 bvector1_reg_0__5_ ( .D(n23253), .CK(clk), .Q(n18951), .QN(n28043) );
  DFF_X2 bvector1_reg_0__4_ ( .D(n23252), .CK(clk), .Q(n18914), .QN(n28042) );
  DFF_X2 bvector0_reg_7__15_ ( .D(n23302), .CK(clk), .QN(n27925) );
  DFF_X2 bvector0_reg_7__14_ ( .D(n23301), .CK(clk), .QN(n27924) );
  DFF_X2 bvector0_reg_7__13_ ( .D(n23300), .CK(clk), .QN(n27923) );
  DFF_X2 bvector0_reg_7__12_ ( .D(n23299), .CK(clk), .QN(n27922) );
  DFF_X2 bvector0_reg_7__11_ ( .D(n23298), .CK(clk), .QN(n27921) );
  DFF_X2 bvector0_reg_7__10_ ( .D(n23297), .CK(clk), .QN(n27920) );
  DFF_X2 bvector0_reg_7__9_ ( .D(n23296), .CK(clk), .QN(n27919) );
  DFF_X2 bvector0_reg_7__8_ ( .D(n23295), .CK(clk), .QN(n27918) );
  DFF_X2 bvector0_reg_7__7_ ( .D(n23294), .CK(clk), .QN(n27917) );
  DFF_X2 bvector0_reg_7__6_ ( .D(n23293), .CK(clk), .QN(n27916) );
  DFF_X2 bvector0_reg_7__5_ ( .D(n23292), .CK(clk), .QN(n27915) );
  DFF_X2 bvector0_reg_7__4_ ( .D(n23291), .CK(clk), .QN(n27914) );
  DFF_X2 bvector0_reg_6__15_ ( .D(n23318), .CK(clk), .QN(n27941) );
  DFF_X2 bvector0_reg_6__14_ ( .D(n23317), .CK(clk), .QN(n27940) );
  DFF_X2 bvector0_reg_6__13_ ( .D(n23316), .CK(clk), .QN(n27939) );
  DFF_X2 bvector0_reg_6__12_ ( .D(n23315), .CK(clk), .QN(n27938) );
  DFF_X2 bvector0_reg_6__11_ ( .D(n23314), .CK(clk), .QN(n27937) );
  DFF_X2 bvector0_reg_6__10_ ( .D(n23313), .CK(clk), .QN(n27936) );
  DFF_X2 bvector0_reg_6__9_ ( .D(n23312), .CK(clk), .QN(n27935) );
  DFF_X2 bvector0_reg_6__8_ ( .D(n23311), .CK(clk), .QN(n27934) );
  DFF_X2 bvector0_reg_6__7_ ( .D(n23310), .CK(clk), .QN(n27933) );
  DFF_X2 bvector0_reg_6__6_ ( .D(n23309), .CK(clk), .QN(n27932) );
  DFF_X2 bvector0_reg_6__5_ ( .D(n23308), .CK(clk), .QN(n27931) );
  DFF_X2 bvector0_reg_6__4_ ( .D(n23307), .CK(clk), .QN(n27930) );
  DFF_X2 bvector0_reg_1__15_ ( .D(n23334), .CK(clk), .QN(n27957) );
  DFF_X2 bvector0_reg_1__14_ ( .D(n23333), .CK(clk), .QN(n27956) );
  DFF_X2 bvector0_reg_1__13_ ( .D(n23332), .CK(clk), .QN(n27955) );
  DFF_X2 z_reg_0__15_ ( .D(n25774), .CK(clk), .QN(n19539) );
  DFF_X2 z_reg_60__15_ ( .D(n25100), .CK(clk), .Q(n26171) );
  DFF_X2 z_reg_59__15_ ( .D(n25384), .CK(clk), .Q(n26159) );
  DFF_X2 z_reg_54__15_ ( .D(n25383), .CK(clk), .Q(n26185), .QN(n19517) );
  DFF_X2 z_reg_51__15_ ( .D(n25382), .CK(clk), .Q(n26188), .QN(n19516) );
  DFF_X2 z_reg_12__15_ ( .D(n25381), .CK(clk), .Q(n26172), .QN(n19545) );
  DFF_X2 z_reg_9__15_ ( .D(n25380), .CK(clk), .Q(n26176), .QN(n19544) );
  DFF_X2 z_reg_4__15_ ( .D(n25379), .CK(clk), .Q(n26145), .QN(n19541) );
  DFF_X2 z_reg_1__15_ ( .D(n25378), .CK(clk), .Q(n26149), .QN(n19540) );
  DFF_X2 z_reg_22__15_ ( .D(n25377), .CK(clk), .Q(n26184), .QN(n19533) );
  DFF_X2 z_reg_19__15_ ( .D(n25376), .CK(clk), .Q(n26187), .QN(n19532) );
  DFF_X2 z_reg_36__15_ ( .D(n25375), .CK(clk), .Q(n26144), .QN(n19525) );
  DFF_X2 z_reg_33__15_ ( .D(n25374), .CK(clk), .Q(n26148), .QN(n19524) );
  DFF_X2 z_reg_30__15_ ( .D(n25096), .CK(clk), .Q(n26156) );
  DFF_X2 z_reg_27__15_ ( .D(n25373), .CK(clk), .Q(n26158) );
  DFF_X2 z_reg_44__15_ ( .D(n25099), .CK(clk), .Q(n26170) );
  DFF_X2 z_reg_41__15_ ( .D(n25372), .CK(clk), .Q(n26175) );
  DFF_X2 z_reg_58__15_ ( .D(n25098), .CK(clk), .Q(n26161) );
  DFF_X2 z_reg_61__15_ ( .D(n25371), .CK(clk), .Q(n26179), .QN(n19522) );
  DFF_X2 z_reg_55__15_ ( .D(n25370), .CK(clk), .Q(n26191) );
  DFF_X2 z_reg_26__15_ ( .D(n25085), .CK(clk), .Q(n26160) );
  DFF_X2 z_reg_18__15_ ( .D(n25369), .CK(clk), .Q(n26189), .QN(n19531) );
  DFF_X2 z_reg_32__15_ ( .D(n25368), .CK(clk), .Q(n26150), .QN(n19523) );
  DFF_X2 z_reg_40__15_ ( .D(n25084), .CK(clk), .Q(n26177) );
  DFF_X2 z_reg_45__15_ ( .D(n25367), .CK(clk), .Q(n26173), .QN(n19530) );
  DFF_X2 z_reg_37__15_ ( .D(n25366), .CK(clk), .Q(n26146) );
  DFF_X2 z_reg_31__15_ ( .D(n25365), .CK(clk), .Q(n26157), .QN(n19538) );
  DFF_X2 z_reg_23__15_ ( .D(n25364), .CK(clk), .Q(n26186) );
  DFF_X2 z_reg_13__15_ ( .D(n25363), .CK(clk), .Q(n26174) );
  DFF_X2 z_reg_5__15_ ( .D(n25362), .CK(clk), .Q(n26147) );
  DFF_X2 z_reg_8__15_ ( .D(n25082), .CK(clk), .Q(n26178) );
  DFF_X2 z_reg_50__15_ ( .D(n25080), .CK(clk), .Q(n26190) );
  DFF_X2 z_reg_9__3_ ( .D(n20735), .CK(clk), .QN(n20324) );
  DFF_X2 z_reg_9__2_ ( .D(n20734), .CK(clk), .QN(n20389) );
  DFF_X2 z_reg_9__1_ ( .D(n20733), .CK(clk), .QN(n20454) );
  DFF_X2 z_reg_9__0_ ( .D(n20732), .CK(clk), .QN(n20520) );
  DFF_X2 z_reg_12__3_ ( .D(n20959), .CK(clk), .QN(n20325) );
  DFF_X2 z_reg_12__2_ ( .D(n20958), .CK(clk), .QN(n20390) );
  DFF_X2 z_reg_12__1_ ( .D(n20957), .CK(clk), .QN(n20455) );
  DFF_X2 z_reg_12__0_ ( .D(n20956), .CK(clk), .QN(n20521) );
  DFF_X2 z_reg_60__3_ ( .D(n20991), .CK(clk), .Q(n28428), .QN(n20301) );
  DFF_X2 z_reg_60__2_ ( .D(n20990), .CK(clk), .Q(n28416), .QN(n20366) );
  DFF_X2 z_reg_60__1_ ( .D(n20989), .CK(clk), .Q(n28404), .QN(n20431) );
  DFF_X2 z_reg_60__0_ ( .D(n20988), .CK(clk), .Q(n28392), .QN(n20497) );
  DFF_X2 z_reg_59__3_ ( .D(n20767), .CK(clk), .Q(n28569), .QN(n20300) );
  DFF_X2 z_reg_59__2_ ( .D(n20766), .CK(clk), .Q(n28554), .QN(n20365) );
  DFF_X2 z_reg_59__1_ ( .D(n20765), .CK(clk), .Q(n28539), .QN(n20430) );
  DFF_X2 z_reg_59__0_ ( .D(n20764), .CK(clk), .Q(n28524), .QN(n20496) );
  DFF_X2 z_reg_44__3_ ( .D(n21055), .CK(clk), .Q(n28425), .QN(n20309) );
  DFF_X2 z_reg_44__2_ ( .D(n21054), .CK(clk), .Q(n28413), .QN(n20374) );
  DFF_X2 z_reg_44__1_ ( .D(n21053), .CK(clk), .Q(n28401), .QN(n20439) );
  DFF_X2 z_reg_44__0_ ( .D(n21052), .CK(clk), .Q(n28389), .QN(n20505) );
  DFF_X2 z_reg_41__3_ ( .D(n20831), .CK(clk), .Q(n28426), .QN(n20308) );
  DFF_X2 z_reg_41__2_ ( .D(n20830), .CK(clk), .Q(n28414), .QN(n20373) );
  DFF_X2 z_reg_41__1_ ( .D(n20829), .CK(clk), .Q(n28402), .QN(n20438) );
  DFF_X2 z_reg_41__0_ ( .D(n20828), .CK(clk), .Q(n28390), .QN(n20504) );
  DFF_X2 z_reg_30__3_ ( .D(n21023), .CK(clk), .Q(n28566), .QN(n20317) );
  DFF_X2 z_reg_30__2_ ( .D(n21022), .CK(clk), .Q(n28551), .QN(n20382) );
  DFF_X2 z_reg_30__1_ ( .D(n21021), .CK(clk), .Q(n28536), .QN(n20447) );
  DFF_X2 z_reg_30__0_ ( .D(n21020), .CK(clk), .Q(n28521), .QN(n20513) );
  DFF_X2 z_reg_27__3_ ( .D(n20799), .CK(clk), .Q(n28567), .QN(n20316) );
  DFF_X2 z_reg_27__2_ ( .D(n20798), .CK(clk), .Q(n28552), .QN(n20381) );
  DFF_X2 z_reg_27__1_ ( .D(n20797), .CK(clk), .Q(n28537), .QN(n20446) );
  DFF_X2 z_reg_27__0_ ( .D(n20796), .CK(clk), .Q(n28522), .QN(n20512) );
  DFF_X2 flag_z_reg ( .D(n23443), .CK(clk), .Q(n26137), .QN(n22426) );
  DFF_X2 z_reg_58__3_ ( .D(n20639), .CK(clk), .Q(n28570), .QN(n20299) );
  DFF_X2 z_reg_58__2_ ( .D(n20638), .CK(clk), .Q(n28555), .QN(n20364) );
  DFF_X2 z_reg_58__1_ ( .D(n20637), .CK(clk), .Q(n28540), .QN(n20429) );
  DFF_X2 z_reg_58__0_ ( .D(n20636), .CK(clk), .Q(n28525), .QN(n20495) );
  DFF_X2 startdesign_reg ( .D(n24818), .CK(clk), .Q(n26135), .QN(n22381) );
  DFF_X2 flag_a_reg ( .D(n21149), .CK(clk), .QN(n16374) );
  DFF_X2 z_reg_40__3_ ( .D(n20703), .CK(clk), .Q(n28427), .QN(n20307) );
  DFF_X2 z_reg_40__2_ ( .D(n20702), .CK(clk), .Q(n28415), .QN(n20372) );
  DFF_X2 z_reg_40__1_ ( .D(n20701), .CK(clk), .Q(n28403), .QN(n20437) );
  DFF_X2 z_reg_40__0_ ( .D(n20700), .CK(clk), .Q(n28391), .QN(n20503) );
  DFF_X2 z_reg_26__3_ ( .D(n20671), .CK(clk), .Q(n28568), .QN(n20315) );
  DFF_X2 z_reg_26__2_ ( .D(n20670), .CK(clk), .Q(n28553), .QN(n20380) );
  DFF_X2 z_reg_26__1_ ( .D(n20669), .CK(clk), .Q(n28538), .QN(n20445) );
  DFF_X2 z_reg_26__0_ ( .D(n20668), .CK(clk), .Q(n28523), .QN(n20511) );
  DFF_X2 z_start_reg ( .D(n23451), .CK(clk), .QN(n22399) );
  DFF_X2 z_reg_61__0_ ( .D(n20572), .CK(clk), .QN(n20498) );
  DFF_X2 z_reg_8__3_ ( .D(n20607), .CK(clk), .Q(n28430), .QN(n20323) );
  DFF_X2 z_reg_8__2_ ( .D(n20606), .CK(clk), .Q(n28418), .QN(n20388) );
  DFF_X2 z_reg_8__1_ ( .D(n20605), .CK(clk), .Q(n28406), .QN(n20453) );
  DFF_X2 z_reg_8__0_ ( .D(n20604), .CK(clk), .Q(n28394), .QN(n20519) );
  DFF_X2 z_reg_45__3_ ( .D(n20927), .CK(clk), .QN(n20310) );
  DFF_X2 z_reg_45__2_ ( .D(n20926), .CK(clk), .QN(n20375) );
  DFF_X2 z_reg_45__1_ ( .D(n20925), .CK(clk), .QN(n20440) );
  DFF_X2 z_reg_45__0_ ( .D(n20924), .CK(clk), .QN(n20506) );
  DFF_X2 z_reg_31__3_ ( .D(n20895), .CK(clk), .QN(n20318) );
  DFF_X2 z_reg_31__2_ ( .D(n20894), .CK(clk), .QN(n20383) );
  DFF_X2 z_reg_31__1_ ( .D(n20893), .CK(clk), .QN(n20448) );
  DFF_X2 z_reg_31__0_ ( .D(n20892), .CK(clk), .QN(n20514) );
  DFF_X2 z_reg_13__3_ ( .D(n20863), .CK(clk), .Q(n28429), .QN(n20326) );
  DFF_X2 z_reg_13__2_ ( .D(n20862), .CK(clk), .Q(n28417), .QN(n20391) );
  DFF_X2 z_reg_13__1_ ( .D(n20861), .CK(clk), .Q(n28405), .QN(n20456) );
  DFF_X2 z_reg_13__0_ ( .D(n20860), .CK(clk), .Q(n28393), .QN(n20522) );
  DFF_X2 z_reg_55__14_ ( .D(n20602), .CK(clk), .Q(n28378), .QN(n19583) );
  DFF_X2 z_reg_60__14_ ( .D(n21002), .CK(clk), .Q(n28507), .QN(n19586) );
  DFF_X2 z_reg_60__13_ ( .D(n21001), .CK(clk), .Q(n28500), .QN(n19651) );
  DFF_X2 z_reg_60__12_ ( .D(n21000), .CK(clk), .Q(n28493), .QN(n19716) );
  DFF_X2 z_reg_60__11_ ( .D(n20999), .CK(clk), .Q(n28486), .QN(n19781) );
  DFF_X2 z_reg_60__10_ ( .D(n20998), .CK(clk), .Q(n28479), .QN(n19846) );
  DFF_X2 z_reg_60__9_ ( .D(n20997), .CK(clk), .Q(n28472), .QN(n19911) );
  DFF_X2 z_reg_60__8_ ( .D(n20996), .CK(clk), .Q(n28465), .QN(n19976) );
  DFF_X2 z_reg_60__7_ ( .D(n20995), .CK(clk), .Q(n28458), .QN(n20041) );
  DFF_X2 z_reg_60__6_ ( .D(n20994), .CK(clk), .Q(n28451), .QN(n20106) );
  DFF_X2 z_reg_60__5_ ( .D(n20993), .CK(clk), .Q(n28444), .QN(n20171) );
  DFF_X2 z_reg_60__4_ ( .D(n20992), .CK(clk), .Q(n28437), .QN(n20236) );
  DFF_X2 z_reg_59__14_ ( .D(n20778), .CK(clk), .Q(n28691), .QN(n19585) );
  DFF_X2 z_reg_59__13_ ( .D(n20777), .CK(clk), .Q(n28680), .QN(n19650) );
  DFF_X2 z_reg_59__12_ ( .D(n20776), .CK(clk), .Q(n28669), .QN(n19715) );
  DFF_X2 z_reg_59__11_ ( .D(n20775), .CK(clk), .Q(n28658), .QN(n19780) );
  DFF_X2 z_reg_59__10_ ( .D(n20774), .CK(clk), .Q(n28647), .QN(n19845) );
  DFF_X2 z_reg_59__9_ ( .D(n20773), .CK(clk), .Q(n28636), .QN(n19910) );
  DFF_X2 z_reg_59__8_ ( .D(n20772), .CK(clk), .Q(n28625), .QN(n19975) );
  DFF_X2 z_reg_59__7_ ( .D(n20771), .CK(clk), .Q(n28614), .QN(n20040) );
  DFF_X2 z_reg_59__6_ ( .D(n20770), .CK(clk), .Q(n28603), .QN(n20105) );
  DFF_X2 z_reg_59__5_ ( .D(n20769), .CK(clk), .Q(n28592), .QN(n20170) );
  DFF_X2 z_reg_59__4_ ( .D(n20768), .CK(clk), .Q(n28581), .QN(n20235) );
  DFF_X2 z_reg_54__14_ ( .D(n21018), .CK(clk), .QN(n19582) );
  DFF_X2 z_reg_54__13_ ( .D(n21017), .CK(clk), .QN(n19647) );
  DFF_X2 z_reg_54__12_ ( .D(n21016), .CK(clk), .QN(n19712) );
  DFF_X2 z_reg_54__11_ ( .D(n21015), .CK(clk), .QN(n19777) );
  DFF_X2 z_reg_54__10_ ( .D(n21014), .CK(clk), .QN(n19842) );
  DFF_X2 z_reg_54__9_ ( .D(n21013), .CK(clk), .QN(n19907) );
  DFF_X2 z_reg_54__8_ ( .D(n21012), .CK(clk), .QN(n19972) );
  DFF_X2 z_reg_54__7_ ( .D(n21011), .CK(clk), .QN(n20037) );
  DFF_X2 sendz_count_reg_0_ ( .D(n23439), .CK(clk), .Q(add_283_A_0_), .QN(
        n22419) );
  DFF_X2 sendz_count_reg_5_ ( .D(n23434), .CK(clk), .Q(add_283_A_5_), .QN(
        n22414) );
  DFF_X2 sendz_count_reg_4_ ( .D(n26297), .CK(clk), .Q(add_283_A_4_), .QN(
        n22415) );
  DFF_X2 sendz_count_reg_3_ ( .D(n26298), .CK(clk), .Q(add_283_A_3_), .QN(
        n22416) );
  DFF_X2 sendz_count_reg_2_ ( .D(n26299), .CK(clk), .Q(add_283_A_2_), .QN(
        n22417) );
  DFF_X2 sendz_count_reg_1_ ( .D(n26300), .CK(clk), .Q(add_283_A_1_), .QN(
        n22418) );
  DFF_X2 bitselect1_reg_1_ ( .D(n23522), .CK(clk), .Q(add_180_A_1_), .QN(
        n22393) );
  DFF_X2 count_m_reg_6_ ( .D(n21160), .CK(clk), .Q(add_1445_B_6_), .QN(n25775)
         );
  DFF_X2 count_m_reg_5_ ( .D(n21159), .CK(clk), .Q(add_1445_B_5_), .QN(n22408)
         );
  DFF_X2 count_m_reg_4_ ( .D(n21158), .CK(clk), .Q(add_1445_B_4_), .QN(n22409)
         );
  DFF_X2 count_m_reg_3_ ( .D(n21157), .CK(clk), .Q(add_1445_B_3_), .QN(n22410)
         );
  DFF_X2 count_m_reg_2_ ( .D(n21156), .CK(clk), .Q(add_1445_B_2_), .QN(n22411)
         );
  DFF_X2 count_m_reg_1_ ( .D(n21155), .CK(clk), .Q(add_1445_B_1_), .QN(n22412)
         );
  DFF_X2 bitselect1_reg_0_ ( .D(n23523), .CK(clk), .Q(add_180_A_0_), .QN(
        n22394) );
  DFF_X2 count_m_reg_0_ ( .D(n23442), .CK(clk), .Q(add_1445_B_0_), .QN(n22413)
         );
  DFF_X2 bitselect1_reg_2_ ( .D(n23521), .CK(clk), .Q(add_180_A_2_), .QN(
        n22392) );
  DFF_X2 count_m_reg_7_ ( .D(n21161), .CK(clk), .Q(add_1445_B_7_), .QN(n18744)
         );
  DFF_X2 count_m_reg_9_ ( .D(n23441), .CK(clk), .Q(add_1445_B_9_), .QN(n22407)
         );
  DFF_X2 bitselect1_reg_3_ ( .D(n23520), .CK(clk), .Q(add_180_A_3_), .QN(
        n22391) );
  DFF_X2 mac_z_reg_15_ ( .D(n20540), .CK(clk), .Q(n651), .QN(n19547) );
  DFF_X2 mac_z_reg_14_ ( .D(n20541), .CK(clk), .Q(n650), .QN(n19612) );
  DFF_X2 mac_z_reg_13_ ( .D(n20542), .CK(clk), .Q(n649), .QN(n19677) );
  DFF_X2 mac_z_reg_12_ ( .D(n20543), .CK(clk), .Q(n648), .QN(n19742) );
  DFF_X2 mac_z_reg_11_ ( .D(n20544), .CK(clk), .Q(n647), .QN(n19807) );
  DFF_X2 mac_z_reg_10_ ( .D(n20545), .CK(clk), .Q(n646), .QN(n19872) );
  DFF_X2 count_m_reg_8_ ( .D(n21162), .CK(clk), .Q(add_1445_B_8_), .QN(n18745)
         );
  DFF_X2 mac_b_reg_15_ ( .D(n23088), .CK(clk), .QN(n25961) );
  DFF_X2 mac_b_reg_14_ ( .D(n23089), .CK(clk), .QN(n25963) );
  DFF_X2 mac_b_reg_13_ ( .D(n23090), .CK(clk), .QN(n25965) );
  DFF_X2 mac_b_reg_12_ ( .D(n23091), .CK(clk), .QN(n25967) );
  DFF_X2 mac_a0_reg_15_ ( .D(n23467), .CK(clk), .Q(n4967), .QN(n18187) );
  DFF_X2 mac_a0_reg_14_ ( .D(n23466), .CK(clk), .Q(n4966), .QN(n18224) );
  DFF_X2 mac_a0_reg_13_ ( .D(n23465), .CK(clk), .Q(n4965), .QN(n18261) );
  DFF_X2 mac_a0_reg_12_ ( .D(n23464), .CK(clk), .Q(n4964), .QN(n18298) );
  DFF_X2 mac_a3_reg_15_ ( .D(n23515), .CK(clk), .Q(n4919), .QN(n16411) );
  DFF_X2 mac_a3_reg_14_ ( .D(n23514), .CK(clk), .Q(n4918), .QN(n16448) );
  DFF_X2 mac_a3_reg_13_ ( .D(n23513), .CK(clk), .Q(n4917), .QN(n16485) );
  DFF_X2 mac_a3_reg_12_ ( .D(n23512), .CK(clk), .Q(n4916), .QN(n16522) );
  DFF_X2 mac_a3_reg_11_ ( .D(n23511), .CK(clk), .Q(n4915), .QN(n16559) );
  DFF_X2 mac_a2_reg_15_ ( .D(n23499), .CK(clk), .Q(n4935), .QN(n17003) );
  DFF_X2 mac_a2_reg_14_ ( .D(n23498), .CK(clk), .Q(n4934), .QN(n17040) );
  DFF_X2 mac_a2_reg_13_ ( .D(n23497), .CK(clk), .Q(n4933), .QN(n17077) );
  DFF_X2 mac_a2_reg_12_ ( .D(n23496), .CK(clk), .Q(n4932), .QN(n17114) );
  DFF_X2 mac_a1_reg_15_ ( .D(n23483), .CK(clk), .Q(n4951), .QN(n17595) );
  DFF_X2 mac_a1_reg_14_ ( .D(n23482), .CK(clk), .Q(n4950), .QN(n17632) );
  DFF_X2 mac_a1_reg_13_ ( .D(n23481), .CK(clk), .Q(n4949), .QN(n17669) );
  DFF_X2 mac_a1_reg_12_ ( .D(n23480), .CK(clk), .Q(n4948), .QN(n17706) );
  DFF_X2 mac_b_reg_11_ ( .D(n23092), .CK(clk), .QN(n25969) );
  DFF_X2 mac_b_reg_10_ ( .D(n23093), .CK(clk), .QN(n25971) );
  DFF_X2 mac_b_reg_9_ ( .D(n23094), .CK(clk), .QN(n25973) );
  DFF_X2 mac_a1_reg_9_ ( .D(n23477), .CK(clk), .Q(n4945), .QN(n17817) );
  DFF_X2 mac_a1_reg_8_ ( .D(n23476), .CK(clk), .Q(n4944), .QN(n17854) );
  DFF_X2 mac_a1_reg_7_ ( .D(n23475), .CK(clk), .Q(n4943), .QN(n17891) );
  DFF_X2 mac_a1_reg_6_ ( .D(n23474), .CK(clk), .Q(n4942), .QN(n17928) );
  DFF_X2 mac_a1_reg_5_ ( .D(n23473), .CK(clk), .Q(n4941), .QN(n17965) );
  DFF_X2 mac_a1_reg_4_ ( .D(n23472), .CK(clk), .Q(n4940), .QN(n18002) );
  DFF_X2 mac_a1_reg_3_ ( .D(n23471), .CK(clk), .Q(n4939), .QN(n18039) );
  DFF_X2 mac_a1_reg_2_ ( .D(n23470), .CK(clk), .Q(n4938), .QN(n18076) );
  DFF_X2 mac_a1_reg_1_ ( .D(n23469), .CK(clk), .Q(n4937), .QN(n18113) );
  DFF_X2 mac_a1_reg_0_ ( .D(n23468), .CK(clk), .Q(n4936), .QN(n18150) );
  DFF_X2 mac_a0_reg_11_ ( .D(n23463), .CK(clk), .Q(n4963), .QN(n18335) );
  DFF_X2 mac_a0_reg_10_ ( .D(n23462), .CK(clk), .Q(n4962), .QN(n18372) );
  DFF_X2 mac_a0_reg_9_ ( .D(n23461), .CK(clk), .Q(n4961), .QN(n18409) );
  DFF_X2 mac_a0_reg_8_ ( .D(n23460), .CK(clk), .Q(n4960), .QN(n18446) );
  DFF_X2 mac_a0_reg_7_ ( .D(n23459), .CK(clk), .Q(n4959), .QN(n18483) );
  DFF_X2 mac_b_reg_5_ ( .D(n23098), .CK(clk), .QN(n18977) );
  SDFF_X2 mac_b_reg_7_ ( .D(1'b1), .SI(1'b0), .SE(n26012), .CK(clk), .QN(
        n25976) );
  DFF_X1 mac_z_reg_0_ ( .D(n20555), .CK(clk), .Q(n636), .QN(n20523) );
  DFF_X2 mac_b_reg_8_ ( .D(n23095), .CK(clk), .QN(n19088) );
  INV_X8 U10540 ( .A(n25976), .ZN(n25975) );
  INV_X4 U10541 ( .A(n20197), .ZN(n25766) );
  INV_X4 U10542 ( .A(n19088), .ZN(n25974) );
  INV_X4 U10543 ( .A(n20327), .ZN(n25764) );
  INV_X4 U10544 ( .A(n16707), .ZN(n25751) );
  INV_X4 U10545 ( .A(n18940), .ZN(n25741) );
  INV_X8 U10546 ( .A(n18977), .ZN(n25978) );
  INV_X8 U10547 ( .A(n19014), .ZN(n25977) );
  INV_X4 U10548 ( .A(n25973), .ZN(n25972) );
  INV_X4 U10549 ( .A(n25967), .ZN(n25966) );
  INV_X4 U10550 ( .A(n25965), .ZN(n25964) );
  INV_X4 U10551 ( .A(n25971), .ZN(n25970) );
  INV_X4 U10552 ( .A(n25969), .ZN(n25968) );
  NAND4_X2 U10553 ( .A1(n11435), .A2(n22422), .A3(n22424), .A4(n24891), .ZN(
        n11645) );
  NAND4_X2 U10554 ( .A1(n11435), .A2(n22422), .A3(n22423), .A4(n24868), .ZN(
        n11641) );
  INV_X4 U10555 ( .A(n16818), .ZN(n25762) );
  NAND2_X2 U10556 ( .A1(n12058), .A2(n24865), .ZN(n24834) );
  NAND2_X2 U10557 ( .A1(n12058), .A2(n12140), .ZN(n24835) );
  NAND2_X2 U10558 ( .A1(n12058), .A2(n12145), .ZN(n24836) );
  NAND2_X2 U10559 ( .A1(n12140), .A2(n12057), .ZN(n24837) );
  NAND2_X2 U10560 ( .A1(n12056), .A2(n12057), .ZN(n24838) );
  NAND2_X2 U10561 ( .A1(n12145), .A2(n12057), .ZN(n24839) );
  NAND2_X2 U10562 ( .A1(n12060), .A2(n12140), .ZN(n24840) );
  NAND2_X2 U10563 ( .A1(n12060), .A2(n24865), .ZN(n24841) );
  NAND2_X2 U10564 ( .A1(n12060), .A2(n12145), .ZN(n24842) );
  NAND2_X2 U10565 ( .A1(n12140), .A2(n12062), .ZN(n24843) );
  NAND2_X2 U10566 ( .A1(n12056), .A2(n12062), .ZN(n24844) );
  NAND2_X2 U10567 ( .A1(n12062), .A2(n24865), .ZN(n24845) );
  NAND2_X2 U10568 ( .A1(n12057), .A2(n24865), .ZN(n24846) );
  AND2_X4 U10569 ( .A1(n12813), .A2(n15479), .ZN(n24847) );
  AND2_X4 U10570 ( .A1(n12813), .A2(n15478), .ZN(n24848) );
  AND2_X4 U10571 ( .A1(n12799), .A2(n15479), .ZN(n24849) );
  AND2_X4 U10572 ( .A1(n12799), .A2(n15478), .ZN(n24850) );
  AND2_X4 U10573 ( .A1(n12812), .A2(n15479), .ZN(n24851) );
  AND2_X4 U10574 ( .A1(n27799), .A2(n15480), .ZN(n24852) );
  AND2_X4 U10575 ( .A1(n12811), .A2(n15479), .ZN(n24853) );
  AND2_X4 U10576 ( .A1(n12786), .A2(n15479), .ZN(n24854) );
  AND2_X4 U10577 ( .A1(n12811), .A2(n15480), .ZN(n24855) );
  AND2_X4 U10578 ( .A1(n12788), .A2(n15480), .ZN(n24856) );
  AND2_X4 U10579 ( .A1(n12803), .A2(n15479), .ZN(n24857) );
  AND2_X4 U10580 ( .A1(n27800), .A2(n15479), .ZN(n24858) );
  AND2_X4 U10581 ( .A1(n12788), .A2(n15478), .ZN(n24859) );
  AND2_X4 U10582 ( .A1(n12803), .A2(n15478), .ZN(n24860) );
  AND2_X4 U10583 ( .A1(n27800), .A2(n15477), .ZN(n24861) );
  AND2_X4 U10584 ( .A1(n12811), .A2(n15477), .ZN(n24862) );
  AND2_X4 U10585 ( .A1(n12786), .A2(n15477), .ZN(n24863) );
  NAND2_X2 U10586 ( .A1(n12062), .A2(n12145), .ZN(n24864) );
  AND2_X4 U10587 ( .A1(n24887), .A2(n25253), .ZN(n24865) );
  AND2_X4 U10588 ( .A1(n27799), .A2(n15477), .ZN(n24866) );
  AND2_X4 U10589 ( .A1(n12811), .A2(n15478), .ZN(n24867) );
  NAND2_X2 U10590 ( .A1(n12799), .A2(n15480), .ZN(n24869) );
  NAND2_X2 U10591 ( .A1(n12799), .A2(n15477), .ZN(n24870) );
  NAND2_X2 U10592 ( .A1(n12803), .A2(n15480), .ZN(n24871) );
  NAND2_X2 U10593 ( .A1(n12803), .A2(n15477), .ZN(n24872) );
  NAND2_X2 U10594 ( .A1(n12812), .A2(n15478), .ZN(n24873) );
  NAND2_X2 U10595 ( .A1(n12812), .A2(n15480), .ZN(n24874) );
  NAND2_X2 U10596 ( .A1(n12812), .A2(n15477), .ZN(n24875) );
  NAND2_X2 U10597 ( .A1(n12788), .A2(n15479), .ZN(n24876) );
  NAND2_X2 U10598 ( .A1(n12813), .A2(n15480), .ZN(n24877) );
  NAND2_X2 U10599 ( .A1(n12813), .A2(n15477), .ZN(n24878) );
  NAND2_X2 U10600 ( .A1(n27799), .A2(n15479), .ZN(n24879) );
  NAND2_X2 U10601 ( .A1(n27799), .A2(n15478), .ZN(n24880) );
  NAND2_X2 U10602 ( .A1(n12786), .A2(n15478), .ZN(n24881) );
  NAND2_X2 U10603 ( .A1(n12786), .A2(n15480), .ZN(n24882) );
  NAND2_X2 U10604 ( .A1(n27800), .A2(n15478), .ZN(n24883) );
  NAND2_X2 U10605 ( .A1(n27800), .A2(n15480), .ZN(n24884) );
  AND2_X4 U10606 ( .A1(n12788), .A2(n15477), .ZN(n24885) );
  AND2_X4 U10607 ( .A1(n24892), .A2(n25251), .ZN(n24886) );
  NAND2_X2 U10608 ( .A1(n12058), .A2(n12056), .ZN(n24888) );
  NAND2_X2 U10609 ( .A1(n12060), .A2(n12056), .ZN(n24889) );
  AND2_X4 U10610 ( .A1(n22414), .A2(n22415), .ZN(n24892) );
  AND2_X4 U10611 ( .A1(n19352), .A2(n26343), .ZN(n24893) );
  AND2_X4 U10612 ( .A1(n11809), .A2(n19356), .ZN(n24897) );
  AND2_X4 U10613 ( .A1(n11806), .A2(n19355), .ZN(n24898) );
  AND2_X4 U10614 ( .A1(n24845), .A2(n26190), .ZN(n25080) );
  AND2_X4 U10615 ( .A1(n24845), .A2(n19487), .ZN(n25081) );
  AND2_X4 U10616 ( .A1(n24864), .A2(n26178), .ZN(n25082) );
  AND2_X4 U10617 ( .A1(n24864), .A2(n19507), .ZN(n25083) );
  AND2_X4 U10618 ( .A1(n25943), .A2(n26177), .ZN(n25084) );
  AND2_X4 U10619 ( .A1(n25946), .A2(n26160), .ZN(n25085) );
  AND2_X4 U10620 ( .A1(n25943), .A2(n19491), .ZN(n25086) );
  AND2_X4 U10621 ( .A1(n25943), .A2(n19495), .ZN(n25087) );
  AND2_X4 U10622 ( .A1(n25946), .A2(n19499), .ZN(n25088) );
  AND2_X4 U10623 ( .A1(n25946), .A2(n19503), .ZN(n25089) );
  AND2_X4 U10624 ( .A1(n25934), .A2(n19500), .ZN(n25090) );
  AND2_X4 U10625 ( .A1(n24889), .A2(n19504), .ZN(n25091) );
  AND2_X4 U10626 ( .A1(n25955), .A2(n19486), .ZN(n25092) );
  AND2_X4 U10627 ( .A1(n25955), .A2(n19490), .ZN(n25093) );
  AND2_X4 U10628 ( .A1(n25931), .A2(n19492), .ZN(n25094) );
  AND2_X4 U10629 ( .A1(n25931), .A2(n19496), .ZN(n25095) );
  AND2_X4 U10630 ( .A1(n25913), .A2(n26156), .ZN(n25096) );
  AND2_X4 U10631 ( .A1(n25919), .A2(n19513), .ZN(n25097) );
  AND2_X4 U10632 ( .A1(n24845), .A2(n26161), .ZN(n25098) );
  AND2_X4 U10633 ( .A1(n25910), .A2(n26170), .ZN(n25099) );
  AND2_X4 U10634 ( .A1(n25916), .A2(n26171), .ZN(n25100) );
  AND2_X4 U10635 ( .A1(n24845), .A2(n19483), .ZN(n25101) );
  AND2_X4 U10636 ( .A1(n25928), .A2(n19514), .ZN(n25102) );
  AND2_X4 U10637 ( .A1(n25940), .A2(n19508), .ZN(n25103) );
  AND2_X4 U10638 ( .A1(n22416), .A2(n22417), .ZN(n25247) );
  AND2_X4 U10639 ( .A1(n22391), .A2(add_180_A_1_), .ZN(n25250) );
  AND2_X4 U10640 ( .A1(n22418), .A2(n22419), .ZN(n25251) );
  AND2_X4 U10641 ( .A1(n11815), .A2(n26162), .ZN(n25258) );
  AND2_X4 U10642 ( .A1(n11813), .A2(n26163), .ZN(n25259) );
  AND2_X4 U10643 ( .A1(n11811), .A2(n26164), .ZN(n25260) );
  AND2_X4 U10644 ( .A1(n11803), .A2(n26165), .ZN(n25261) );
  AND2_X4 U10645 ( .A1(n11801), .A2(n26166), .ZN(n25262) );
  AND2_X4 U10646 ( .A1(n24864), .A2(n26151), .ZN(n25361) );
  AND2_X4 U10647 ( .A1(n24839), .A2(n26147), .ZN(n25362) );
  AND2_X4 U10648 ( .A1(n25928), .A2(n26174), .ZN(n25363) );
  AND2_X4 U10649 ( .A1(n24838), .A2(n26186), .ZN(n25364) );
  AND2_X4 U10650 ( .A1(n25925), .A2(n26157), .ZN(n25365) );
  AND2_X4 U10651 ( .A1(n24837), .A2(n26146), .ZN(n25366) );
  AND2_X4 U10652 ( .A1(n25922), .A2(n26173), .ZN(n25367) );
  AND2_X4 U10653 ( .A1(n24843), .A2(n26150), .ZN(n25368) );
  AND2_X4 U10654 ( .A1(n24844), .A2(n26189), .ZN(n25369) );
  AND2_X4 U10655 ( .A1(n25955), .A2(n26191), .ZN(n25370) );
  AND2_X4 U10656 ( .A1(n25955), .A2(n26179), .ZN(n25371) );
  AND2_X4 U10657 ( .A1(n24840), .A2(n26175), .ZN(n25372) );
  AND2_X4 U10658 ( .A1(n25934), .A2(n26158), .ZN(n25373) );
  AND2_X4 U10659 ( .A1(n25931), .A2(n26148), .ZN(n25374) );
  AND2_X4 U10660 ( .A1(n24835), .A2(n26144), .ZN(n25375) );
  AND2_X4 U10661 ( .A1(n25934), .A2(n26187), .ZN(n25376) );
  AND2_X4 U10662 ( .A1(n25913), .A2(n26184), .ZN(n25377) );
  AND2_X4 U10663 ( .A1(n24842), .A2(n26149), .ZN(n25378) );
  AND2_X4 U10664 ( .A1(n24836), .A2(n26145), .ZN(n25379) );
  AND2_X4 U10665 ( .A1(n25940), .A2(n26176), .ZN(n25380) );
  AND2_X4 U10666 ( .A1(n25919), .A2(n26172), .ZN(n25381) );
  AND2_X4 U10667 ( .A1(n24841), .A2(n26188), .ZN(n25382) );
  AND2_X4 U10668 ( .A1(n24834), .A2(n26185), .ZN(n25383) );
  AND2_X4 U10669 ( .A1(n25937), .A2(n26159), .ZN(n25384) );
  AND2_X4 U10670 ( .A1(n25928), .A2(n26180), .ZN(n25385) );
  AND2_X4 U10671 ( .A1(n25925), .A2(n26143), .ZN(n25386) );
  AND2_X4 U10672 ( .A1(n25925), .A2(n26169), .ZN(n25387) );
  AND2_X4 U10673 ( .A1(n25922), .A2(n26183), .ZN(n25388) );
  AND2_X4 U10674 ( .A1(n25922), .A2(n26155), .ZN(n25389) );
  AND2_X4 U10675 ( .A1(n25910), .A2(n26182), .ZN(n25390) );
  AND2_X4 U10676 ( .A1(n25910), .A2(n26154), .ZN(n25391) );
  AND2_X4 U10677 ( .A1(n25913), .A2(n26142), .ZN(n25392) );
  AND2_X4 U10678 ( .A1(n24888), .A2(n26168), .ZN(n25393) );
  AND2_X4 U10679 ( .A1(n25919), .A2(n26181), .ZN(n25394) );
  AND2_X4 U10680 ( .A1(n25940), .A2(n26152), .ZN(n25395) );
  AND2_X4 U10681 ( .A1(n25937), .A2(n26140), .ZN(n25396) );
  AND2_X4 U10682 ( .A1(n24834), .A2(n26141), .ZN(n25397) );
  AND2_X4 U10683 ( .A1(n25937), .A2(n26167), .ZN(n25398) );
  AND2_X4 U10684 ( .A1(n24834), .A2(n26153), .ZN(n25399) );
  INV_X1 U10685 ( .A(n25742), .ZN(n25732) );
  INV_X4 U10688 ( .A(n25735), .ZN(n25736) );
  INV_X4 U10689 ( .A(n20526), .ZN(n25737) );
  INV_X4 U10690 ( .A(n18903), .ZN(n25980) );
  INV_X4 U10691 ( .A(n16966), .ZN(n25752) );
  INV_X4 U10692 ( .A(n20529), .ZN(n25738) );
  INV_X4 U10693 ( .A(n25739), .ZN(n25740) );
  INV_X4 U10694 ( .A(n18940), .ZN(n25979) );
  INV_X2 U10695 ( .A(n25769), .ZN(n25742) );
  INV_X4 U10696 ( .A(n25743), .ZN(n25744) );
  INV_X4 U10697 ( .A(n25745), .ZN(n25746) );
  INV_X2 U10698 ( .A(n20262), .ZN(n25759) );
  INV_X4 U10699 ( .A(n20392), .ZN(n25747) );
  INV_X4 U10700 ( .A(n20528), .ZN(n25748) );
  INV_X4 U10701 ( .A(n25749), .ZN(n25750) );
  INV_X1 U10702 ( .A(n25983), .ZN(n25753) );
  INV_X4 U10703 ( .A(n25753), .ZN(n25754) );
  INV_X4 U10704 ( .A(n25984), .ZN(n25983) );
  INV_X4 U10705 ( .A(n25755), .ZN(n25756) );
  MUX2_X1 U10706 ( .A(n25756), .B(n26133), .S(n25959), .Z(n25986) );
  INV_X2 U10707 ( .A(n20525), .ZN(n25760) );
  INV_X4 U10708 ( .A(n25757), .ZN(n25758) );
  INV_X4 U10709 ( .A(n18866), .ZN(n25761) );
  INV_X4 U10710 ( .A(n25982), .ZN(n25981) );
  MUX2_X1 U10711 ( .A(n25746), .B(n26023), .S(n25907), .Z(n26024) );
  INV_X4 U10712 ( .A(n16929), .ZN(n25763) );
  MUX2_X1 U10713 ( .A(n25744), .B(n25999), .S(n26130), .Z(n26000) );
  INV_X4 U10714 ( .A(n16781), .ZN(n25780) );
  MUX2_X1 U10715 ( .A(n25758), .B(n25991), .S(n26130), .Z(n25992) );
  INV_X4 U10716 ( .A(n20457), .ZN(n25767) );
  MUX2_X1 U10717 ( .A(n25736), .B(n26031), .S(n25907), .Z(n26032) );
  INV_X2 U10718 ( .A(n16855), .ZN(n25765) );
  AOI221_X1 U10719 ( .B1(n19352), .B2(n11647), .C1(n26303), .C2(
        dut__dom__data[15]), .A(n11789), .ZN(n11779) );
  AOI221_X1 U10720 ( .B1(n19360), .B2(n11647), .C1(n26303), .C2(
        dut__dom__data[14]), .A(n11776), .ZN(n11770) );
  AOI221_X1 U10721 ( .B1(n19368), .B2(n11647), .C1(n26303), .C2(
        dut__dom__data[13]), .A(n11767), .ZN(n11761) );
  AOI221_X1 U10722 ( .B1(n19376), .B2(n11647), .C1(n26303), .C2(
        dut__dom__data[12]), .A(n11758), .ZN(n11752) );
  AOI221_X1 U10723 ( .B1(n19384), .B2(n11647), .C1(n26303), .C2(
        dut__dom__data[11]), .A(n11749), .ZN(n11743) );
  AOI221_X1 U10724 ( .B1(n19392), .B2(n11647), .C1(n26303), .C2(
        dut__dom__data[10]), .A(n11740), .ZN(n11734) );
  AOI221_X1 U10725 ( .B1(n19400), .B2(n11647), .C1(n26303), .C2(
        dut__dom__data[9]), .A(n11731), .ZN(n11725) );
  AOI221_X1 U10726 ( .B1(n19408), .B2(n11647), .C1(n26303), .C2(
        dut__dom__data[8]), .A(n11722), .ZN(n11716) );
  AOI221_X1 U10727 ( .B1(n19416), .B2(n11647), .C1(n26303), .C2(
        dut__dom__data[7]), .A(n11713), .ZN(n11707) );
  AOI221_X1 U10728 ( .B1(n19424), .B2(n11647), .C1(n26303), .C2(
        dut__dom__data[6]), .A(n11704), .ZN(n11698) );
  AOI221_X1 U10729 ( .B1(n19432), .B2(n11647), .C1(n26303), .C2(
        dut__dom__data[5]), .A(n11695), .ZN(n11689) );
  AOI221_X1 U10730 ( .B1(n19440), .B2(n11647), .C1(n26303), .C2(
        dut__dom__data[4]), .A(n11686), .ZN(n11680) );
  AOI221_X1 U10731 ( .B1(n19448), .B2(n11647), .C1(n26303), .C2(
        dut__dom__data[3]), .A(n11677), .ZN(n11671) );
  AOI221_X1 U10732 ( .B1(n19456), .B2(n11647), .C1(n26303), .C2(
        dut__dom__data[2]), .A(n11668), .ZN(n11662) );
  AOI221_X1 U10733 ( .B1(n19464), .B2(n11647), .C1(n26303), .C2(
        dut__dom__data[1]), .A(n11659), .ZN(n11653) );
  AOI221_X1 U10734 ( .B1(n19472), .B2(n11647), .C1(n26303), .C2(
        dut__dom__data[0]), .A(n11648), .ZN(n11636) );
  INV_X4 U10735 ( .A(n25961), .ZN(n25960) );
  INV_X4 U10736 ( .A(n25963), .ZN(n25962) );
  INV_X4 U10737 ( .A(n24866), .ZN(n25884) );
  INV_X4 U10738 ( .A(n24866), .ZN(n25883) );
  INV_X4 U10739 ( .A(n24852), .ZN(n25880) );
  INV_X4 U10740 ( .A(n24852), .ZN(n25879) );
  INV_X4 U10741 ( .A(n24879), .ZN(n25886) );
  INV_X4 U10742 ( .A(n24879), .ZN(n25885) );
  INV_X4 U10743 ( .A(n24880), .ZN(n25888) );
  INV_X4 U10744 ( .A(n24880), .ZN(n25887) );
  INV_X4 U10745 ( .A(n25930), .ZN(n25928) );
  INV_X4 U10746 ( .A(n24850), .ZN(n25900) );
  INV_X4 U10747 ( .A(n24850), .ZN(n25899) );
  INV_X4 U10748 ( .A(n24849), .ZN(n25902) );
  INV_X4 U10749 ( .A(n24849), .ZN(n25901) );
  INV_X4 U10750 ( .A(n24853), .ZN(n25844) );
  INV_X4 U10751 ( .A(n24853), .ZN(n25843) );
  INV_X4 U10752 ( .A(n24861), .ZN(n25898) );
  INV_X4 U10753 ( .A(n24861), .ZN(n25897) );
  INV_X4 U10754 ( .A(n24855), .ZN(n25846) );
  INV_X4 U10755 ( .A(n24855), .ZN(n25845) );
  INV_X4 U10756 ( .A(n24867), .ZN(n25847) );
  INV_X4 U10757 ( .A(n24867), .ZN(n25848) );
  INV_X4 U10758 ( .A(n24883), .ZN(n25903) );
  INV_X4 U10759 ( .A(n24869), .ZN(n25839) );
  INV_X4 U10760 ( .A(n24883), .ZN(n25904) );
  INV_X4 U10761 ( .A(n24869), .ZN(n25840) );
  INV_X4 U10762 ( .A(n24870), .ZN(n25842) );
  INV_X4 U10763 ( .A(n24870), .ZN(n25841) );
  INV_X4 U10764 ( .A(n24884), .ZN(n25906) );
  INV_X4 U10765 ( .A(n24884), .ZN(n25905) );
  INV_X4 U10766 ( .A(n24862), .ZN(n25855) );
  INV_X4 U10767 ( .A(n24862), .ZN(n25856) );
  INV_X4 U10768 ( .A(n24858), .ZN(n25890) );
  INV_X4 U10769 ( .A(n24858), .ZN(n25889) );
  INV_X4 U10770 ( .A(n24839), .ZN(n25929) );
  INV_X4 U10771 ( .A(n24839), .ZN(n25930) );
  INV_X4 U10772 ( .A(n25957), .ZN(n25955) );
  INV_X4 U10773 ( .A(n25954), .ZN(n25952) );
  INV_X4 U10774 ( .A(n25942), .ZN(n25940) );
  INV_X4 U10775 ( .A(n25921), .ZN(n25919) );
  INV_X4 U10776 ( .A(n25945), .ZN(n25943) );
  INV_X4 U10777 ( .A(n25933), .ZN(n25931) );
  INV_X4 U10778 ( .A(n25912), .ZN(n25910) );
  INV_X4 U10779 ( .A(n25924), .ZN(n25922) );
  INV_X4 U10780 ( .A(n25939), .ZN(n25937) );
  INV_X4 U10781 ( .A(n25948), .ZN(n25946) );
  INV_X4 U10782 ( .A(n25936), .ZN(n25934) );
  INV_X4 U10783 ( .A(n25915), .ZN(n25913) );
  INV_X4 U10784 ( .A(n25927), .ZN(n25925) );
  INV_X4 U10785 ( .A(n25918), .ZN(n25916) );
  INV_X4 U10786 ( .A(dim__dut__data[12]), .ZN(n25792) );
  INV_X4 U10787 ( .A(dim__dut__data[11]), .ZN(n25797) );
  INV_X4 U10788 ( .A(dim__dut__data[1]), .ZN(n25828) );
  INV_X4 U10789 ( .A(dim__dut__data[15]), .ZN(n25783) );
  INV_X4 U10790 ( .A(dim__dut__data[14]), .ZN(n25786) );
  INV_X4 U10791 ( .A(dim__dut__data[13]), .ZN(n25789) );
  INV_X4 U10792 ( .A(dim__dut__data[12]), .ZN(n25794) );
  INV_X4 U10793 ( .A(dim__dut__data[11]), .ZN(n25799) );
  INV_X4 U10794 ( .A(dim__dut__data[10]), .ZN(n25801) );
  INV_X4 U10795 ( .A(dim__dut__data[9]), .ZN(n25804) );
  INV_X4 U10796 ( .A(dim__dut__data[8]), .ZN(n25807) );
  INV_X4 U10797 ( .A(dim__dut__data[7]), .ZN(n25810) );
  INV_X4 U10798 ( .A(dim__dut__data[6]), .ZN(n25813) );
  INV_X4 U10799 ( .A(dim__dut__data[5]), .ZN(n25816) );
  INV_X4 U10800 ( .A(dim__dut__data[4]), .ZN(n25819) );
  INV_X4 U10801 ( .A(dim__dut__data[3]), .ZN(n25822) );
  INV_X4 U10802 ( .A(dim__dut__data[2]), .ZN(n25825) );
  INV_X4 U10803 ( .A(dim__dut__data[1]), .ZN(n25830) );
  INV_X4 U10804 ( .A(dim__dut__data[0]), .ZN(n25833) );
  INV_X4 U10805 ( .A(dim__dut__data[15]), .ZN(n25784) );
  INV_X4 U10806 ( .A(dim__dut__data[14]), .ZN(n25787) );
  INV_X4 U10807 ( .A(dim__dut__data[13]), .ZN(n25790) );
  INV_X4 U10808 ( .A(dim__dut__data[12]), .ZN(n25795) );
  INV_X4 U10809 ( .A(dim__dut__data[10]), .ZN(n25802) );
  INV_X4 U10810 ( .A(dim__dut__data[9]), .ZN(n25805) );
  INV_X4 U10811 ( .A(dim__dut__data[8]), .ZN(n25808) );
  INV_X4 U10812 ( .A(dim__dut__data[7]), .ZN(n25811) );
  INV_X4 U10813 ( .A(dim__dut__data[6]), .ZN(n25814) );
  INV_X4 U10814 ( .A(dim__dut__data[5]), .ZN(n25817) );
  INV_X4 U10815 ( .A(dim__dut__data[4]), .ZN(n25820) );
  INV_X4 U10816 ( .A(dim__dut__data[3]), .ZN(n25823) );
  INV_X4 U10817 ( .A(dim__dut__data[2]), .ZN(n25826) );
  INV_X4 U10818 ( .A(dim__dut__data[1]), .ZN(n25831) );
  INV_X4 U10819 ( .A(dim__dut__data[0]), .ZN(n25834) );
  INV_X4 U10820 ( .A(dim__dut__data[12]), .ZN(n25791) );
  INV_X4 U10821 ( .A(dim__dut__data[11]), .ZN(n25796) );
  INV_X4 U10822 ( .A(dim__dut__data[1]), .ZN(n25827) );
  INV_X4 U10823 ( .A(dim__dut__data[15]), .ZN(n25782) );
  INV_X4 U10824 ( .A(dim__dut__data[14]), .ZN(n25785) );
  INV_X4 U10825 ( .A(dim__dut__data[13]), .ZN(n25788) );
  INV_X4 U10826 ( .A(dim__dut__data[12]), .ZN(n25793) );
  INV_X4 U10827 ( .A(dim__dut__data[11]), .ZN(n25798) );
  INV_X4 U10828 ( .A(dim__dut__data[10]), .ZN(n25800) );
  INV_X4 U10829 ( .A(dim__dut__data[9]), .ZN(n25803) );
  INV_X4 U10830 ( .A(dim__dut__data[8]), .ZN(n25806) );
  INV_X4 U10831 ( .A(dim__dut__data[7]), .ZN(n25809) );
  INV_X4 U10832 ( .A(dim__dut__data[6]), .ZN(n25812) );
  INV_X4 U10833 ( .A(dim__dut__data[5]), .ZN(n25815) );
  INV_X4 U10834 ( .A(dim__dut__data[4]), .ZN(n25818) );
  INV_X4 U10835 ( .A(dim__dut__data[3]), .ZN(n25821) );
  INV_X4 U10836 ( .A(dim__dut__data[2]), .ZN(n25824) );
  INV_X4 U10837 ( .A(dim__dut__data[1]), .ZN(n25829) );
  INV_X4 U10838 ( .A(dim__dut__data[0]), .ZN(n25832) );
  NAND2_X2 U10839 ( .A1(n27799), .A2(n12791), .ZN(n12210) );
  NAND2_X2 U10840 ( .A1(n27799), .A2(n12790), .ZN(n12226) );
  INV_X4 U10841 ( .A(n25959), .ZN(n25958) );
  INV_X4 U10842 ( .A(n24856), .ZN(n25866) );
  INV_X4 U10843 ( .A(n24856), .ZN(n25865) );
  INV_X4 U10844 ( .A(n24885), .ZN(n25864) );
  INV_X4 U10845 ( .A(n24885), .ZN(n25863) );
  INV_X4 U10846 ( .A(n24859), .ZN(n25862) );
  INV_X4 U10847 ( .A(n24859), .ZN(n25861) );
  INV_X4 U10848 ( .A(n24854), .ZN(n25881) );
  INV_X4 U10849 ( .A(n24854), .ZN(n25882) );
  NAND2_X2 U10850 ( .A1(n27799), .A2(n12787), .ZN(n12201) );
  INV_X4 U10851 ( .A(n25908), .ZN(n25907) );
  INV_X4 U10852 ( .A(n24875), .ZN(n25867) );
  INV_X4 U10853 ( .A(n24881), .ZN(n25893) );
  INV_X4 U10854 ( .A(n24873), .ZN(n25857) );
  INV_X4 U10855 ( .A(n24877), .ZN(n25875) );
  INV_X4 U10856 ( .A(n24871), .ZN(n25849) );
  INV_X4 U10857 ( .A(n24881), .ZN(n25894) );
  INV_X4 U10858 ( .A(n24875), .ZN(n25868) );
  INV_X4 U10859 ( .A(n24873), .ZN(n25858) );
  INV_X4 U10860 ( .A(n24877), .ZN(n25876) );
  INV_X4 U10861 ( .A(n24871), .ZN(n25850) );
  INV_X4 U10862 ( .A(n24878), .ZN(n25878) );
  INV_X4 U10863 ( .A(n24876), .ZN(n25870) );
  INV_X4 U10864 ( .A(n24872), .ZN(n25852) );
  INV_X4 U10865 ( .A(n24876), .ZN(n25869) );
  INV_X4 U10866 ( .A(n24872), .ZN(n25851) );
  INV_X4 U10867 ( .A(n24878), .ZN(n25877) );
  INV_X4 U10868 ( .A(n24882), .ZN(n25896) );
  INV_X4 U10869 ( .A(n24874), .ZN(n25860) );
  INV_X4 U10870 ( .A(n24882), .ZN(n25895) );
  INV_X4 U10871 ( .A(n24874), .ZN(n25859) );
  INV_X4 U10872 ( .A(n24857), .ZN(n25838) );
  INV_X4 U10873 ( .A(n24847), .ZN(n25873) );
  INV_X4 U10874 ( .A(n24857), .ZN(n25837) );
  INV_X4 U10875 ( .A(n24847), .ZN(n25874) );
  INV_X4 U10876 ( .A(n24848), .ZN(n25871) );
  INV_X4 U10877 ( .A(n24860), .ZN(n25835) );
  INV_X4 U10878 ( .A(n24848), .ZN(n25872) );
  INV_X4 U10879 ( .A(n24860), .ZN(n25836) );
  INV_X4 U10880 ( .A(n24863), .ZN(n25891) );
  INV_X4 U10881 ( .A(n24863), .ZN(n25892) );
  INV_X4 U10882 ( .A(n24851), .ZN(n25854) );
  INV_X4 U10883 ( .A(n24851), .ZN(n25853) );
  INV_X4 U10884 ( .A(n11798), .ZN(n26343) );
  INV_X4 U10885 ( .A(n12843), .ZN(n26337) );
  INV_X4 U10886 ( .A(n12892), .ZN(n26328) );
  INV_X4 U10887 ( .A(n12980), .ZN(n26319) );
  INV_X4 U10888 ( .A(n12872), .ZN(n26333) );
  INV_X4 U10889 ( .A(n12853), .ZN(n26334) );
  INV_X4 U10890 ( .A(n12849), .ZN(n26335) );
  INV_X4 U10891 ( .A(n12846), .ZN(n26336) );
  INV_X4 U10892 ( .A(n12948), .ZN(n26324) );
  INV_X4 U10893 ( .A(n12930), .ZN(n26325) );
  INV_X4 U10894 ( .A(n12927), .ZN(n26326) );
  INV_X4 U10895 ( .A(n12910), .ZN(n26327) );
  INV_X4 U10896 ( .A(n12988), .ZN(n26315) );
  INV_X4 U10897 ( .A(n12986), .ZN(n26316) );
  INV_X4 U10898 ( .A(n12984), .ZN(n26317) );
  INV_X4 U10899 ( .A(n12982), .ZN(n26318) );
  INV_X4 U10900 ( .A(n13012), .ZN(n26308) );
  INV_X4 U10901 ( .A(n16300), .ZN(n26464) );
  INV_X4 U10902 ( .A(n16240), .ZN(n26473) );
  INV_X4 U10903 ( .A(n16137), .ZN(n26482) );
  INV_X4 U10904 ( .A(n16078), .ZN(n26491) );
  INV_X4 U10905 ( .A(n16051), .ZN(n26425) );
  INV_X4 U10906 ( .A(n16025), .ZN(n26434) );
  INV_X4 U10907 ( .A(n15999), .ZN(n26443) );
  INV_X4 U10908 ( .A(n15972), .ZN(n26452) );
  INV_X4 U10909 ( .A(n15930), .ZN(n26389) );
  INV_X4 U10910 ( .A(n15888), .ZN(n26398) );
  INV_X4 U10911 ( .A(n15846), .ZN(n26407) );
  INV_X4 U10912 ( .A(n15803), .ZN(n26416) );
  INV_X4 U10913 ( .A(n15743), .ZN(n26353) );
  INV_X4 U10914 ( .A(n15686), .ZN(n26362) );
  INV_X4 U10915 ( .A(n15628), .ZN(n26371) );
  INV_X4 U10916 ( .A(n15569), .ZN(n26380) );
  INV_X4 U10917 ( .A(n13031), .ZN(n26306) );
  INV_X4 U10918 ( .A(n16321), .ZN(n26462) );
  INV_X4 U10919 ( .A(n16261), .ZN(n26471) );
  INV_X4 U10920 ( .A(n16158), .ZN(n26480) );
  INV_X4 U10921 ( .A(n16099), .ZN(n26489) );
  INV_X4 U10922 ( .A(n16055), .ZN(n26423) );
  INV_X4 U10923 ( .A(n16029), .ZN(n26432) );
  INV_X4 U10924 ( .A(n16003), .ZN(n26441) );
  INV_X4 U10925 ( .A(n15976), .ZN(n26450) );
  INV_X4 U10926 ( .A(n15949), .ZN(n26387) );
  INV_X4 U10927 ( .A(n15907), .ZN(n26396) );
  INV_X4 U10928 ( .A(n15865), .ZN(n26405) );
  INV_X4 U10929 ( .A(n15822), .ZN(n26414) );
  INV_X4 U10930 ( .A(n15764), .ZN(n26351) );
  INV_X4 U10931 ( .A(n15707), .ZN(n26360) );
  INV_X4 U10932 ( .A(n15649), .ZN(n26369) );
  INV_X4 U10933 ( .A(n15590), .ZN(n26378) );
  INV_X4 U10934 ( .A(n13029), .ZN(n26307) );
  INV_X4 U10935 ( .A(n16303), .ZN(n26463) );
  INV_X4 U10936 ( .A(n16243), .ZN(n26472) );
  INV_X4 U10937 ( .A(n16140), .ZN(n26481) );
  INV_X4 U10938 ( .A(n16081), .ZN(n26490) );
  INV_X4 U10939 ( .A(n16053), .ZN(n26424) );
  INV_X4 U10940 ( .A(n16027), .ZN(n26433) );
  INV_X4 U10941 ( .A(n16001), .ZN(n26442) );
  INV_X4 U10942 ( .A(n15974), .ZN(n26451) );
  INV_X4 U10943 ( .A(n15947), .ZN(n26388) );
  INV_X4 U10944 ( .A(n15905), .ZN(n26397) );
  INV_X4 U10945 ( .A(n15863), .ZN(n26406) );
  INV_X4 U10946 ( .A(n15820), .ZN(n26415) );
  INV_X4 U10947 ( .A(n15746), .ZN(n26352) );
  INV_X4 U10948 ( .A(n15689), .ZN(n26361) );
  INV_X4 U10949 ( .A(n15631), .ZN(n26370) );
  INV_X4 U10950 ( .A(n15572), .ZN(n26379) );
  INV_X4 U10951 ( .A(n12992), .ZN(n26310) );
  INV_X4 U10952 ( .A(n16118), .ZN(n26484) );
  INV_X4 U10953 ( .A(n16279), .ZN(n26466) );
  INV_X4 U10954 ( .A(n15979), .ZN(n26445) );
  INV_X4 U10955 ( .A(n15825), .ZN(n26409) );
  INV_X4 U10956 ( .A(n15609), .ZN(n26373) );
  INV_X4 U10957 ( .A(n16221), .ZN(n26475) );
  INV_X4 U10958 ( .A(n16031), .ZN(n26427) );
  INV_X4 U10959 ( .A(n15867), .ZN(n26400) );
  INV_X4 U10960 ( .A(n16059), .ZN(n26493) );
  INV_X4 U10961 ( .A(n15909), .ZN(n26391) );
  INV_X4 U10962 ( .A(n16005), .ZN(n26436) );
  INV_X4 U10963 ( .A(n15667), .ZN(n26364) );
  INV_X4 U10964 ( .A(n15952), .ZN(n26454) );
  INV_X4 U10965 ( .A(n15550), .ZN(n26382) );
  INV_X4 U10966 ( .A(n15782), .ZN(n26418) );
  INV_X4 U10967 ( .A(n11430), .ZN(n26355) );
  INV_X4 U10968 ( .A(n15741), .ZN(n26354) );
  INV_X4 U10969 ( .A(n13009), .ZN(n26309) );
  INV_X4 U10970 ( .A(n16296), .ZN(n26465) );
  INV_X4 U10971 ( .A(n16238), .ZN(n26474) );
  INV_X4 U10972 ( .A(n16135), .ZN(n26483) );
  INV_X4 U10973 ( .A(n16076), .ZN(n26492) );
  INV_X4 U10974 ( .A(n16034), .ZN(n26426) );
  INV_X4 U10975 ( .A(n16008), .ZN(n26435) );
  INV_X4 U10976 ( .A(n15982), .ZN(n26444) );
  INV_X4 U10977 ( .A(n15955), .ZN(n26453) );
  INV_X4 U10978 ( .A(n15912), .ZN(n26390) );
  INV_X4 U10979 ( .A(n15870), .ZN(n26399) );
  INV_X4 U10980 ( .A(n15828), .ZN(n26408) );
  INV_X4 U10981 ( .A(n15785), .ZN(n26417) );
  INV_X4 U10982 ( .A(n15684), .ZN(n26363) );
  INV_X4 U10983 ( .A(n15626), .ZN(n26372) );
  INV_X4 U10984 ( .A(n15567), .ZN(n26381) );
  INV_X4 U10985 ( .A(n11452), .ZN(n26341) );
  INV_X4 U10986 ( .A(n11455), .ZN(n26340) );
  INV_X4 U10987 ( .A(n11457), .ZN(n26339) );
  INV_X4 U10988 ( .A(n11459), .ZN(n26338) );
  INV_X4 U10989 ( .A(n11461), .ZN(n26332) );
  INV_X4 U10990 ( .A(n11464), .ZN(n26331) );
  INV_X4 U10991 ( .A(n11466), .ZN(n26330) );
  INV_X4 U10992 ( .A(n11468), .ZN(n26329) );
  INV_X4 U10993 ( .A(n11470), .ZN(n26323) );
  INV_X4 U10994 ( .A(n11473), .ZN(n26322) );
  INV_X4 U10995 ( .A(n11475), .ZN(n26321) );
  INV_X4 U10996 ( .A(n11477), .ZN(n26320) );
  INV_X4 U10997 ( .A(n11428), .ZN(n26356) );
  INV_X4 U10998 ( .A(n11425), .ZN(n26357) );
  INV_X4 U10999 ( .A(n11402), .ZN(n26359) );
  INV_X4 U11000 ( .A(n11479), .ZN(n26314) );
  INV_X4 U11001 ( .A(n11482), .ZN(n26313) );
  INV_X4 U11002 ( .A(n11484), .ZN(n26312) );
  INV_X4 U11003 ( .A(n11486), .ZN(n26311) );
  INV_X4 U11004 ( .A(n11505), .ZN(n26468) );
  INV_X4 U11005 ( .A(n11541), .ZN(n26429) );
  INV_X4 U11006 ( .A(n11577), .ZN(n26393) );
  INV_X4 U11007 ( .A(n11500), .ZN(n26470) );
  INV_X4 U11008 ( .A(n11536), .ZN(n26431) );
  INV_X4 U11009 ( .A(n11572), .ZN(n26395) );
  INV_X4 U11010 ( .A(n11503), .ZN(n26469) );
  INV_X4 U11011 ( .A(n11539), .ZN(n26430) );
  INV_X4 U11012 ( .A(n11575), .ZN(n26394) );
  INV_X4 U11013 ( .A(n11507), .ZN(n26467) );
  INV_X4 U11014 ( .A(n11543), .ZN(n26428) );
  INV_X4 U11015 ( .A(n11579), .ZN(n26392) );
  INV_X4 U11016 ( .A(n11514), .ZN(n26477) );
  INV_X4 U11017 ( .A(n11523), .ZN(n26486) );
  INV_X4 U11018 ( .A(n11532), .ZN(n26495) );
  INV_X4 U11019 ( .A(n11550), .ZN(n26438) );
  INV_X4 U11020 ( .A(n11559), .ZN(n26447) );
  INV_X4 U11021 ( .A(n11568), .ZN(n26456) );
  INV_X4 U11022 ( .A(n11586), .ZN(n26402) );
  INV_X4 U11023 ( .A(n11595), .ZN(n26411) );
  INV_X4 U11024 ( .A(n11604), .ZN(n26420) );
  INV_X4 U11025 ( .A(n11613), .ZN(n26366) );
  INV_X4 U11026 ( .A(n11622), .ZN(n26375) );
  INV_X4 U11027 ( .A(n11631), .ZN(n26384) );
  INV_X4 U11028 ( .A(n11509), .ZN(n26479) );
  INV_X4 U11029 ( .A(n11518), .ZN(n26488) );
  INV_X4 U11030 ( .A(n11527), .ZN(n26497) );
  INV_X4 U11031 ( .A(n11545), .ZN(n26440) );
  INV_X4 U11032 ( .A(n11554), .ZN(n26449) );
  INV_X4 U11033 ( .A(n11563), .ZN(n26458) );
  INV_X4 U11034 ( .A(n11581), .ZN(n26404) );
  INV_X4 U11035 ( .A(n11590), .ZN(n26413) );
  INV_X4 U11036 ( .A(n11599), .ZN(n26422) );
  INV_X4 U11037 ( .A(n11608), .ZN(n26368) );
  INV_X4 U11038 ( .A(n11617), .ZN(n26377) );
  INV_X4 U11039 ( .A(n11626), .ZN(n26386) );
  INV_X4 U11040 ( .A(n11512), .ZN(n26478) );
  INV_X4 U11041 ( .A(n11521), .ZN(n26487) );
  INV_X4 U11042 ( .A(n11530), .ZN(n26496) );
  INV_X4 U11043 ( .A(n11548), .ZN(n26439) );
  INV_X4 U11044 ( .A(n11557), .ZN(n26448) );
  INV_X4 U11045 ( .A(n11566), .ZN(n26457) );
  INV_X4 U11046 ( .A(n11584), .ZN(n26403) );
  INV_X4 U11047 ( .A(n11593), .ZN(n26412) );
  INV_X4 U11048 ( .A(n11602), .ZN(n26421) );
  INV_X4 U11049 ( .A(n11611), .ZN(n26367) );
  INV_X4 U11050 ( .A(n11620), .ZN(n26376) );
  INV_X4 U11051 ( .A(n11629), .ZN(n26385) );
  INV_X4 U11052 ( .A(n11516), .ZN(n26476) );
  INV_X4 U11053 ( .A(n11525), .ZN(n26485) );
  INV_X4 U11054 ( .A(n11534), .ZN(n26494) );
  INV_X4 U11055 ( .A(n11552), .ZN(n26437) );
  INV_X4 U11056 ( .A(n11561), .ZN(n26446) );
  INV_X4 U11057 ( .A(n11570), .ZN(n26455) );
  INV_X4 U11058 ( .A(n11588), .ZN(n26401) );
  INV_X4 U11059 ( .A(n11597), .ZN(n26410) );
  INV_X4 U11060 ( .A(n11606), .ZN(n26419) );
  INV_X4 U11061 ( .A(n11615), .ZN(n26365) );
  INV_X4 U11062 ( .A(n11624), .ZN(n26374) );
  INV_X4 U11063 ( .A(n11633), .ZN(n26383) );
  INV_X4 U11064 ( .A(n11422), .ZN(n26358) );
  INV_X4 U11065 ( .A(n24845), .ZN(n25950) );
  INV_X4 U11066 ( .A(n24841), .ZN(n25938) );
  INV_X4 U11067 ( .A(n24834), .ZN(n25917) );
  INV_X4 U11068 ( .A(n24844), .ZN(n25947) );
  INV_X4 U11069 ( .A(n24889), .ZN(n25935) );
  INV_X4 U11070 ( .A(n24888), .ZN(n25914) );
  INV_X4 U11071 ( .A(n24838), .ZN(n25926) );
  INV_X4 U11072 ( .A(n24864), .ZN(n25953) );
  INV_X4 U11073 ( .A(n24842), .ZN(n25941) );
  INV_X4 U11074 ( .A(n24836), .ZN(n25920) );
  INV_X4 U11075 ( .A(n24843), .ZN(n25944) );
  INV_X4 U11076 ( .A(n24840), .ZN(n25932) );
  INV_X4 U11077 ( .A(n24835), .ZN(n25911) );
  INV_X4 U11078 ( .A(n24837), .ZN(n25923) );
  INV_X4 U11079 ( .A(n24846), .ZN(n25956) );
  INV_X4 U11080 ( .A(n24864), .ZN(n25954) );
  INV_X4 U11081 ( .A(n24842), .ZN(n25942) );
  INV_X4 U11082 ( .A(n24836), .ZN(n25921) );
  INV_X4 U11083 ( .A(n24843), .ZN(n25945) );
  INV_X4 U11084 ( .A(n24840), .ZN(n25933) );
  INV_X4 U11085 ( .A(n24835), .ZN(n25912) );
  INV_X4 U11086 ( .A(n24837), .ZN(n25924) );
  INV_X4 U11087 ( .A(n24845), .ZN(n25951) );
  INV_X4 U11088 ( .A(n24841), .ZN(n25939) );
  INV_X4 U11089 ( .A(n24834), .ZN(n25918) );
  INV_X4 U11090 ( .A(n24844), .ZN(n25948) );
  INV_X4 U11091 ( .A(n24889), .ZN(n25936) );
  INV_X4 U11092 ( .A(n24888), .ZN(n25915) );
  INV_X4 U11093 ( .A(n24838), .ZN(n25927) );
  INV_X4 U11094 ( .A(n24846), .ZN(n25957) );
  INV_X4 U11095 ( .A(n25951), .ZN(n25949) );
  NAND2_X2 U11096 ( .A1(n12811), .A2(n12789), .ZN(n12215) );
  NAND4_X2 U11097 ( .A1(n12814), .A2(n12815), .A3(n12816), .A4(n12817), .ZN(
        n12787) );
  NAND4_X2 U11098 ( .A1(n12825), .A2(n12826), .A3(n12827), .A4(n12828), .ZN(
        n12791) );
  NAND4_X2 U11099 ( .A1(n12838), .A2(n12839), .A3(n12840), .A4(n12841), .ZN(
        n12790) );
  INV_X4 U11100 ( .A(n12972), .ZN(n26500) );
  NAND4_X2 U11101 ( .A1(n12829), .A2(n12830), .A3(n12831), .A4(n12832), .ZN(
        n12789) );
  NAND2_X2 U11102 ( .A1(n27800), .A2(n12787), .ZN(n12175) );
  INV_X4 U11103 ( .A(n12971), .ZN(n26508) );
  NAND4_X2 U11104 ( .A1(n12816), .A2(n12828), .A3(n12832), .A4(n12841), .ZN(
        n15479) );
  NAND4_X2 U11105 ( .A1(n12814), .A2(n12825), .A3(n12829), .A4(n12838), .ZN(
        n15477) );
  NAND4_X2 U11106 ( .A1(n12817), .A2(n12827), .A3(n12831), .A4(n12840), .ZN(
        n15478) );
  AOI21_X2 U11107 ( .B1(n15780), .B2(n26518), .A(n26460), .ZN(n16179) );
  NAND4_X2 U11108 ( .A1(n12815), .A2(n12826), .A3(n12830), .A4(n12839), .ZN(
        n15480) );
  INV_X4 U11109 ( .A(n11878), .ZN(n26139) );
  INV_X4 U11110 ( .A(n11811), .ZN(n26346) );
  INV_X4 U11111 ( .A(n25909), .ZN(n25908) );
  NAND2_X2 U11112 ( .A1(n12799), .A2(n12787), .ZN(n12180) );
  INV_X4 U11113 ( .A(n11283), .ZN(n25959) );
  NAND2_X2 U11114 ( .A1(n12799), .A2(n12791), .ZN(n12183) );
  NAND2_X2 U11115 ( .A1(n27800), .A2(n12790), .ZN(n12182) );
  NAND2_X2 U11116 ( .A1(n12811), .A2(n12787), .ZN(n12200) );
  NOR2_X2 U11117 ( .A1(n26303), .A2(n26305), .ZN(n11647) );
  NOR2_X2 U11118 ( .A1(n13043), .A2(n25958), .ZN(n11798) );
  NAND2_X2 U11119 ( .A1(n12844), .A2(n11419), .ZN(n11430) );
  NAND2_X2 U11120 ( .A1(n11419), .A2(n26502), .ZN(n11402) );
  NAND2_X2 U11121 ( .A1(n11453), .A2(n25781), .ZN(n11455) );
  NAND2_X2 U11122 ( .A1(n11453), .A2(n12844), .ZN(n12843) );
  NAND2_X2 U11123 ( .A1(n11462), .A2(n25781), .ZN(n11464) );
  NAND2_X2 U11124 ( .A1(n11462), .A2(n12844), .ZN(n12892) );
  NAND2_X2 U11125 ( .A1(n11471), .A2(n25781), .ZN(n11473) );
  NAND2_X2 U11126 ( .A1(n11471), .A2(n12844), .ZN(n12980) );
  NAND2_X2 U11127 ( .A1(n11480), .A2(n25781), .ZN(n11482) );
  NAND2_X2 U11128 ( .A1(n11480), .A2(n12844), .ZN(n12992) );
  NAND2_X2 U11129 ( .A1(n11501), .A2(n25781), .ZN(n11503) );
  NAND2_X2 U11130 ( .A1(n11519), .A2(n12844), .ZN(n16118) );
  NAND2_X2 U11131 ( .A1(n11510), .A2(n25781), .ZN(n11512) );
  NAND2_X2 U11132 ( .A1(n11519), .A2(n25781), .ZN(n11521) );
  NAND2_X2 U11133 ( .A1(n11528), .A2(n25781), .ZN(n11530) );
  NAND2_X2 U11134 ( .A1(n11537), .A2(n25781), .ZN(n11539) );
  NAND2_X2 U11135 ( .A1(n11546), .A2(n25781), .ZN(n11548) );
  NAND2_X2 U11136 ( .A1(n11555), .A2(n25781), .ZN(n11557) );
  NAND2_X2 U11137 ( .A1(n11564), .A2(n25781), .ZN(n11566) );
  NAND2_X2 U11138 ( .A1(n11573), .A2(n25781), .ZN(n11575) );
  NAND2_X2 U11139 ( .A1(n11582), .A2(n25781), .ZN(n11584) );
  NAND2_X2 U11140 ( .A1(n11591), .A2(n25781), .ZN(n11593) );
  NAND2_X2 U11141 ( .A1(n11600), .A2(n25781), .ZN(n11602) );
  NAND2_X2 U11142 ( .A1(n11609), .A2(n25781), .ZN(n11611) );
  NAND2_X2 U11143 ( .A1(n11618), .A2(n25781), .ZN(n11620) );
  NAND2_X2 U11144 ( .A1(n11627), .A2(n25781), .ZN(n11629) );
  NAND2_X2 U11145 ( .A1(n11555), .A2(n12844), .ZN(n15979) );
  NAND2_X2 U11146 ( .A1(n11591), .A2(n12844), .ZN(n15825) );
  NAND2_X2 U11147 ( .A1(n11618), .A2(n12844), .ZN(n15609) );
  NAND2_X2 U11148 ( .A1(n11510), .A2(n12844), .ZN(n16221) );
  NAND2_X2 U11149 ( .A1(n11546), .A2(n12844), .ZN(n16005) );
  NAND2_X2 U11150 ( .A1(n11582), .A2(n12844), .ZN(n15867) );
  NAND2_X2 U11151 ( .A1(n11609), .A2(n12844), .ZN(n15667) );
  NAND2_X2 U11152 ( .A1(n11537), .A2(n12844), .ZN(n16031) );
  NAND2_X2 U11153 ( .A1(n11564), .A2(n12844), .ZN(n15952) );
  NAND2_X2 U11154 ( .A1(n11501), .A2(n12844), .ZN(n16279) );
  NAND2_X2 U11155 ( .A1(n11528), .A2(n12844), .ZN(n16059) );
  NAND2_X2 U11156 ( .A1(n11627), .A2(n12844), .ZN(n15550) );
  NAND2_X2 U11157 ( .A1(n11573), .A2(n12844), .ZN(n15909) );
  NAND2_X2 U11158 ( .A1(n11600), .A2(n12844), .ZN(n15782) );
  NAND2_X2 U11159 ( .A1(n26506), .A2(n11453), .ZN(n12872) );
  NAND2_X2 U11160 ( .A1(n26510), .A2(n11453), .ZN(n12853) );
  NAND2_X2 U11161 ( .A1(n11453), .A2(n26502), .ZN(n11452) );
  NAND2_X2 U11162 ( .A1(n11453), .A2(n26500), .ZN(n11457) );
  NAND2_X2 U11163 ( .A1(n11453), .A2(n26509), .ZN(n11459) );
  NAND2_X2 U11164 ( .A1(n26508), .A2(n11453), .ZN(n12849) );
  NAND2_X2 U11165 ( .A1(n12847), .A2(n11453), .ZN(n12846) );
  NAND2_X2 U11166 ( .A1(n26506), .A2(n11462), .ZN(n12948) );
  NAND2_X2 U11167 ( .A1(n26510), .A2(n11462), .ZN(n12930) );
  NAND2_X2 U11168 ( .A1(n11462), .A2(n26502), .ZN(n11461) );
  NAND2_X2 U11169 ( .A1(n11462), .A2(n26500), .ZN(n11466) );
  NAND2_X2 U11170 ( .A1(n11462), .A2(n26509), .ZN(n11468) );
  NAND2_X2 U11171 ( .A1(n26508), .A2(n11462), .ZN(n12927) );
  NAND2_X2 U11172 ( .A1(n12847), .A2(n11462), .ZN(n12910) );
  NAND2_X2 U11173 ( .A1(n26506), .A2(n11471), .ZN(n12988) );
  NAND2_X2 U11174 ( .A1(n26510), .A2(n11471), .ZN(n12986) );
  NAND2_X2 U11175 ( .A1(n11471), .A2(n26502), .ZN(n11470) );
  NAND2_X2 U11176 ( .A1(n11471), .A2(n26500), .ZN(n11475) );
  NAND2_X2 U11177 ( .A1(n11471), .A2(n26509), .ZN(n11477) );
  NAND2_X2 U11178 ( .A1(n26508), .A2(n11471), .ZN(n12984) );
  NAND2_X2 U11179 ( .A1(n12847), .A2(n11471), .ZN(n12982) );
  NAND2_X2 U11180 ( .A1(n26506), .A2(n11480), .ZN(n13031) );
  NAND2_X2 U11181 ( .A1(n26510), .A2(n11480), .ZN(n13029) );
  NAND2_X2 U11182 ( .A1(n11480), .A2(n26502), .ZN(n11479) );
  NAND2_X2 U11183 ( .A1(n11480), .A2(n26500), .ZN(n11484) );
  NAND2_X2 U11184 ( .A1(n11480), .A2(n26509), .ZN(n11486) );
  NAND2_X2 U11185 ( .A1(n26508), .A2(n11480), .ZN(n13012) );
  NAND2_X2 U11186 ( .A1(n12847), .A2(n11480), .ZN(n13009) );
  NAND2_X2 U11187 ( .A1(n11501), .A2(n26500), .ZN(n11505) );
  NAND2_X2 U11188 ( .A1(n11510), .A2(n26500), .ZN(n11514) );
  NAND2_X2 U11189 ( .A1(n11519), .A2(n26500), .ZN(n11523) );
  NAND2_X2 U11190 ( .A1(n11528), .A2(n26500), .ZN(n11532) );
  NAND2_X2 U11191 ( .A1(n11537), .A2(n26500), .ZN(n11541) );
  NAND2_X2 U11192 ( .A1(n11546), .A2(n26500), .ZN(n11550) );
  NAND2_X2 U11193 ( .A1(n11555), .A2(n26500), .ZN(n11559) );
  NAND2_X2 U11194 ( .A1(n11564), .A2(n26500), .ZN(n11568) );
  NAND2_X2 U11195 ( .A1(n11573), .A2(n26500), .ZN(n11577) );
  NAND2_X2 U11196 ( .A1(n11582), .A2(n26500), .ZN(n11586) );
  NAND2_X2 U11197 ( .A1(n11591), .A2(n26500), .ZN(n11595) );
  NAND2_X2 U11198 ( .A1(n11600), .A2(n26500), .ZN(n11604) );
  NAND2_X2 U11199 ( .A1(n26500), .A2(n11419), .ZN(n11425) );
  NAND2_X2 U11200 ( .A1(n11609), .A2(n26500), .ZN(n11613) );
  NAND2_X2 U11201 ( .A1(n11618), .A2(n26500), .ZN(n11622) );
  NAND2_X2 U11202 ( .A1(n11627), .A2(n26500), .ZN(n11631) );
  NAND2_X2 U11203 ( .A1(n12847), .A2(n11501), .ZN(n16296) );
  NAND2_X2 U11204 ( .A1(n12847), .A2(n11510), .ZN(n16238) );
  NAND2_X2 U11205 ( .A1(n12847), .A2(n11519), .ZN(n16135) );
  NAND2_X2 U11206 ( .A1(n12847), .A2(n11528), .ZN(n16076) );
  NAND2_X2 U11207 ( .A1(n12847), .A2(n11537), .ZN(n16034) );
  NAND2_X2 U11208 ( .A1(n12847), .A2(n11546), .ZN(n16008) );
  NAND2_X2 U11209 ( .A1(n12847), .A2(n11555), .ZN(n15982) );
  NAND2_X2 U11210 ( .A1(n12847), .A2(n11564), .ZN(n15955) );
  NAND2_X2 U11211 ( .A1(n12847), .A2(n11573), .ZN(n15912) );
  NAND2_X2 U11212 ( .A1(n12847), .A2(n11582), .ZN(n15870) );
  NAND2_X2 U11213 ( .A1(n12847), .A2(n11591), .ZN(n15828) );
  NAND2_X2 U11214 ( .A1(n12847), .A2(n11600), .ZN(n15785) );
  NAND2_X2 U11215 ( .A1(n12847), .A2(n11419), .ZN(n15741) );
  NAND2_X2 U11216 ( .A1(n12847), .A2(n11609), .ZN(n15684) );
  NAND2_X2 U11217 ( .A1(n12847), .A2(n11618), .ZN(n15626) );
  NAND2_X2 U11218 ( .A1(n12847), .A2(n11627), .ZN(n15567) );
  NAND2_X2 U11219 ( .A1(n11501), .A2(n26502), .ZN(n11500) );
  NAND2_X2 U11220 ( .A1(n11510), .A2(n26502), .ZN(n11509) );
  NAND2_X2 U11221 ( .A1(n11519), .A2(n26502), .ZN(n11518) );
  NAND2_X2 U11222 ( .A1(n11528), .A2(n26502), .ZN(n11527) );
  NAND2_X2 U11223 ( .A1(n11537), .A2(n26502), .ZN(n11536) );
  NAND2_X2 U11224 ( .A1(n11546), .A2(n26502), .ZN(n11545) );
  NAND2_X2 U11225 ( .A1(n11555), .A2(n26502), .ZN(n11554) );
  NAND2_X2 U11226 ( .A1(n11564), .A2(n26502), .ZN(n11563) );
  NAND2_X2 U11227 ( .A1(n11573), .A2(n26502), .ZN(n11572) );
  NAND2_X2 U11228 ( .A1(n11582), .A2(n26502), .ZN(n11581) );
  NAND2_X2 U11229 ( .A1(n11591), .A2(n26502), .ZN(n11590) );
  NAND2_X2 U11230 ( .A1(n11600), .A2(n26502), .ZN(n11599) );
  NAND2_X2 U11231 ( .A1(n11609), .A2(n26502), .ZN(n11608) );
  NAND2_X2 U11232 ( .A1(n11618), .A2(n26502), .ZN(n11617) );
  NAND2_X2 U11233 ( .A1(n11627), .A2(n26502), .ZN(n11626) );
  NAND2_X2 U11234 ( .A1(n26506), .A2(n11501), .ZN(n16321) );
  NAND2_X2 U11235 ( .A1(n26506), .A2(n11510), .ZN(n16261) );
  NAND2_X2 U11236 ( .A1(n26506), .A2(n11519), .ZN(n16158) );
  NAND2_X2 U11237 ( .A1(n26506), .A2(n11528), .ZN(n16099) );
  NAND2_X2 U11238 ( .A1(n26506), .A2(n11537), .ZN(n16055) );
  NAND2_X2 U11239 ( .A1(n26506), .A2(n11546), .ZN(n16029) );
  NAND2_X2 U11240 ( .A1(n26506), .A2(n11555), .ZN(n16003) );
  NAND2_X2 U11241 ( .A1(n26506), .A2(n11564), .ZN(n15976) );
  NAND2_X2 U11242 ( .A1(n26506), .A2(n11573), .ZN(n15949) );
  NAND2_X2 U11243 ( .A1(n26506), .A2(n11582), .ZN(n15907) );
  NAND2_X2 U11244 ( .A1(n26506), .A2(n11591), .ZN(n15865) );
  NAND2_X2 U11245 ( .A1(n26506), .A2(n11600), .ZN(n15822) );
  NAND2_X2 U11246 ( .A1(n26506), .A2(n11419), .ZN(n15764) );
  NAND2_X2 U11247 ( .A1(n26506), .A2(n11609), .ZN(n15707) );
  NAND2_X2 U11248 ( .A1(n26506), .A2(n11618), .ZN(n15649) );
  NAND2_X2 U11249 ( .A1(n26506), .A2(n11627), .ZN(n15590) );
  NAND2_X2 U11250 ( .A1(n26510), .A2(n11501), .ZN(n16303) );
  NAND2_X2 U11251 ( .A1(n26510), .A2(n11510), .ZN(n16243) );
  NAND2_X2 U11252 ( .A1(n26510), .A2(n11519), .ZN(n16140) );
  NAND2_X2 U11253 ( .A1(n26510), .A2(n11528), .ZN(n16081) );
  NAND2_X2 U11254 ( .A1(n26510), .A2(n11537), .ZN(n16053) );
  NAND2_X2 U11255 ( .A1(n26510), .A2(n11546), .ZN(n16027) );
  NAND2_X2 U11256 ( .A1(n26510), .A2(n11555), .ZN(n16001) );
  NAND2_X2 U11257 ( .A1(n26510), .A2(n11564), .ZN(n15974) );
  NAND2_X2 U11258 ( .A1(n26510), .A2(n11573), .ZN(n15947) );
  NAND2_X2 U11259 ( .A1(n26510), .A2(n11582), .ZN(n15905) );
  NAND2_X2 U11260 ( .A1(n26510), .A2(n11591), .ZN(n15863) );
  NAND2_X2 U11261 ( .A1(n26510), .A2(n11600), .ZN(n15820) );
  NAND2_X2 U11262 ( .A1(n26510), .A2(n11419), .ZN(n15746) );
  NAND2_X2 U11263 ( .A1(n26510), .A2(n11609), .ZN(n15689) );
  NAND2_X2 U11264 ( .A1(n26510), .A2(n11618), .ZN(n15631) );
  NAND2_X2 U11265 ( .A1(n26510), .A2(n11627), .ZN(n15572) );
  NAND2_X2 U11266 ( .A1(n25781), .A2(n11419), .ZN(n11422) );
  NAND2_X2 U11267 ( .A1(n11501), .A2(n26509), .ZN(n11507) );
  NAND2_X2 U11268 ( .A1(n11510), .A2(n26509), .ZN(n11516) );
  NAND2_X2 U11269 ( .A1(n11519), .A2(n26509), .ZN(n11525) );
  NAND2_X2 U11270 ( .A1(n11528), .A2(n26509), .ZN(n11534) );
  NAND2_X2 U11271 ( .A1(n11537), .A2(n26509), .ZN(n11543) );
  NAND2_X2 U11272 ( .A1(n11546), .A2(n26509), .ZN(n11552) );
  NAND2_X2 U11273 ( .A1(n11555), .A2(n26509), .ZN(n11561) );
  NAND2_X2 U11274 ( .A1(n11564), .A2(n26509), .ZN(n11570) );
  NAND2_X2 U11275 ( .A1(n11573), .A2(n26509), .ZN(n11579) );
  NAND2_X2 U11276 ( .A1(n11582), .A2(n26509), .ZN(n11588) );
  NAND2_X2 U11277 ( .A1(n11591), .A2(n26509), .ZN(n11597) );
  NAND2_X2 U11278 ( .A1(n11600), .A2(n26509), .ZN(n11606) );
  NAND2_X2 U11279 ( .A1(n26509), .A2(n11419), .ZN(n11428) );
  NAND2_X2 U11280 ( .A1(n11609), .A2(n26509), .ZN(n11615) );
  NAND2_X2 U11281 ( .A1(n11618), .A2(n26509), .ZN(n11624) );
  NAND2_X2 U11282 ( .A1(n11627), .A2(n26509), .ZN(n11633) );
  NAND2_X2 U11283 ( .A1(n26508), .A2(n11501), .ZN(n16300) );
  NAND2_X2 U11284 ( .A1(n26508), .A2(n11510), .ZN(n16240) );
  NAND2_X2 U11285 ( .A1(n26508), .A2(n11519), .ZN(n16137) );
  NAND2_X2 U11286 ( .A1(n26508), .A2(n11528), .ZN(n16078) );
  NAND2_X2 U11287 ( .A1(n26508), .A2(n11537), .ZN(n16051) );
  NAND2_X2 U11288 ( .A1(n26508), .A2(n11546), .ZN(n16025) );
  NAND2_X2 U11289 ( .A1(n26508), .A2(n11555), .ZN(n15999) );
  NAND2_X2 U11290 ( .A1(n26508), .A2(n11564), .ZN(n15972) );
  NAND2_X2 U11291 ( .A1(n26508), .A2(n11573), .ZN(n15930) );
  NAND2_X2 U11292 ( .A1(n26508), .A2(n11582), .ZN(n15888) );
  NAND2_X2 U11293 ( .A1(n26508), .A2(n11591), .ZN(n15846) );
  NAND2_X2 U11294 ( .A1(n26508), .A2(n11600), .ZN(n15803) );
  NAND2_X2 U11295 ( .A1(n26508), .A2(n11419), .ZN(n15743) );
  NAND2_X2 U11296 ( .A1(n26508), .A2(n11609), .ZN(n15686) );
  NAND2_X2 U11297 ( .A1(n26508), .A2(n11618), .ZN(n15628) );
  NAND2_X2 U11298 ( .A1(n26508), .A2(n11627), .ZN(n15569) );
  INV_X4 U11299 ( .A(n11801), .ZN(n26349) );
  NOR4_X2 U11300 ( .A1(add_180_A_3_), .A2(add_180_A_2_), .A3(add_180_A_1_), 
        .A4(add_180_A_0_), .ZN(n12799) );
  NAND2_X2 U11301 ( .A1(n12788), .A2(n12791), .ZN(n12216) );
  OAI222_X2 U11302 ( .A1(n11641), .A2(n28820), .B1(n11643), .B2(n28821), .C1(
        n11645), .C2(n28819), .ZN(n11781) );
  OAI222_X2 U11303 ( .A1(n11641), .A2(n28815), .B1(n11643), .B2(n28816), .C1(
        n11645), .C2(n28814), .ZN(n11772) );
  OAI222_X2 U11304 ( .A1(n11641), .A2(n28807), .B1(n11643), .B2(n28808), .C1(
        n11645), .C2(n28806), .ZN(n11763) );
  OAI222_X2 U11305 ( .A1(n11641), .A2(n28799), .B1(n11643), .B2(n28800), .C1(
        n11645), .C2(n28798), .ZN(n11754) );
  OAI222_X2 U11306 ( .A1(n11641), .A2(n28791), .B1(n11643), .B2(n28792), .C1(
        n11645), .C2(n28790), .ZN(n11745) );
  OAI222_X2 U11307 ( .A1(n11641), .A2(n28783), .B1(n11643), .B2(n28784), .C1(
        n11645), .C2(n28782), .ZN(n11736) );
  OAI222_X2 U11308 ( .A1(n11641), .A2(n28775), .B1(n11643), .B2(n28776), .C1(
        n11645), .C2(n28774), .ZN(n11727) );
  OAI222_X2 U11309 ( .A1(n11641), .A2(n28767), .B1(n11643), .B2(n28768), .C1(
        n11645), .C2(n28766), .ZN(n11718) );
  OAI222_X2 U11310 ( .A1(n11641), .A2(n28759), .B1(n11643), .B2(n28760), .C1(
        n11645), .C2(n28758), .ZN(n11709) );
  OAI222_X2 U11311 ( .A1(n11641), .A2(n28751), .B1(n11643), .B2(n28752), .C1(
        n11645), .C2(n28750), .ZN(n11700) );
  OAI222_X2 U11312 ( .A1(n11641), .A2(n28743), .B1(n11643), .B2(n28744), .C1(
        n11645), .C2(n28742), .ZN(n11691) );
  OAI222_X2 U11313 ( .A1(n11641), .A2(n28735), .B1(n11643), .B2(n28736), .C1(
        n11645), .C2(n28734), .ZN(n11682) );
  OAI222_X2 U11314 ( .A1(n11641), .A2(n28727), .B1(n11643), .B2(n28728), .C1(
        n11645), .C2(n28726), .ZN(n11673) );
  OAI222_X2 U11315 ( .A1(n11641), .A2(n28719), .B1(n11643), .B2(n28720), .C1(
        n11645), .C2(n28718), .ZN(n11664) );
  OAI222_X2 U11316 ( .A1(n11641), .A2(n28711), .B1(n11643), .B2(n28712), .C1(
        n11645), .C2(n28710), .ZN(n11655) );
  OAI222_X2 U11317 ( .A1(n11641), .A2(n28703), .B1(n11643), .B2(n28704), .C1(
        n11645), .C2(n28702), .ZN(n11640) );
  INV_X4 U11318 ( .A(n16205), .ZN(n26502) );
  NAND2_X2 U11319 ( .A1(n11225), .A2(n25247), .ZN(n10178) );
  NAND2_X2 U11320 ( .A1(n11225), .A2(n11196), .ZN(n10170) );
  NAND2_X2 U11321 ( .A1(n11245), .A2(n11200), .ZN(n10156) );
  NAND2_X2 U11322 ( .A1(n11245), .A2(n11195), .ZN(n10163) );
  NAND2_X2 U11323 ( .A1(n11196), .A2(n11266), .ZN(n10189) );
  NAND2_X2 U11324 ( .A1(n11195), .A2(n11266), .ZN(n10196) );
  NAND2_X2 U11325 ( .A1(n11276), .A2(n11200), .ZN(n10203) );
  NAND2_X2 U11326 ( .A1(n11276), .A2(n11195), .ZN(n10210) );
  NAND2_X2 U11327 ( .A1(n12803), .A2(n12791), .ZN(n12188) );
  NAND2_X2 U11328 ( .A1(n12813), .A2(n12791), .ZN(n12208) );
  NAND2_X2 U11329 ( .A1(n12813), .A2(n12790), .ZN(n12224) );
  NAND2_X2 U11330 ( .A1(n11221), .A2(n11200), .ZN(n10172) );
  NAND2_X2 U11331 ( .A1(n11227), .A2(n11195), .ZN(n10180) );
  NAND2_X2 U11332 ( .A1(n11244), .A2(n11200), .ZN(n10158) );
  NAND2_X2 U11333 ( .A1(n11244), .A2(n11195), .ZN(n10165) );
  NAND2_X2 U11334 ( .A1(n11196), .A2(n11265), .ZN(n10191) );
  NAND2_X2 U11335 ( .A1(n11195), .A2(n11265), .ZN(n10198) );
  NAND2_X2 U11336 ( .A1(n11275), .A2(n11200), .ZN(n10205) );
  NAND2_X2 U11337 ( .A1(n11275), .A2(n11195), .ZN(n10212) );
  NAND2_X2 U11338 ( .A1(n12803), .A2(n12787), .ZN(n12190) );
  NAND2_X2 U11339 ( .A1(n11226), .A2(n25247), .ZN(n10133) );
  NAND2_X2 U11340 ( .A1(n11194), .A2(n25247), .ZN(n10147) );
  NAND2_X2 U11341 ( .A1(n24886), .A2(n25247), .ZN(n10102) );
  NAND2_X2 U11342 ( .A1(n11226), .A2(n11195), .ZN(n10140) );
  NAND2_X2 U11343 ( .A1(n11221), .A2(n11195), .ZN(n10126) );
  NAND2_X2 U11344 ( .A1(n11194), .A2(n11195), .ZN(n10095) );
  NAND2_X2 U11345 ( .A1(n24886), .A2(n11195), .ZN(n10109) );
  NAND2_X2 U11346 ( .A1(n24886), .A2(n11200), .ZN(n10115) );
  INV_X4 U11347 ( .A(n16208), .ZN(n26506) );
  NAND2_X2 U11348 ( .A1(n11231), .A2(n25247), .ZN(n10141) );
  NAND2_X2 U11349 ( .A1(n11220), .A2(n25247), .ZN(n10127) );
  NAND2_X2 U11350 ( .A1(n11192), .A2(n25247), .ZN(n10096) );
  NAND2_X2 U11351 ( .A1(n11207), .A2(n25247), .ZN(n10110) );
  NAND2_X2 U11352 ( .A1(n11207), .A2(n11196), .ZN(n10116) );
  NAND2_X2 U11353 ( .A1(n12786), .A2(n12790), .ZN(n12176) );
  NAND2_X2 U11354 ( .A1(n11225), .A2(n11200), .ZN(n10134) );
  NAND2_X2 U11355 ( .A1(n11231), .A2(n11200), .ZN(n10148) );
  NAND2_X2 U11356 ( .A1(n11192), .A2(n11200), .ZN(n10103) );
  NAND2_X2 U11357 ( .A1(n11634), .A2(n25958), .ZN(n11441) );
  INV_X4 U11358 ( .A(n11435), .ZN(n26303) );
  NOR3_X2 U11359 ( .A1(n24833), .A2(n25400), .A3(n16298), .ZN(n12847) );
  OAI21_X2 U11360 ( .B1(n25104), .B2(n26283), .A(n13091), .ZN(n13086) );
  OAI21_X2 U11361 ( .B1(add_180_A_1_), .B2(n26285), .A(n15545), .ZN(n15541) );
  OAI21_X2 U11362 ( .B1(n26293), .B2(n24868), .A(n16364), .ZN(n16361) );
  NAND2_X2 U11363 ( .A1(n11283), .A2(n12977), .ZN(n11437) );
  OAI21_X2 U11364 ( .B1(n12978), .B2(n11490), .A(n11794), .ZN(n12977) );
  INV_X4 U11365 ( .A(n11815), .ZN(n26344) );
  INV_X4 U11366 ( .A(n11634), .ZN(n26293) );
  NAND2_X2 U11368 ( .A1(n12788), .A2(n12790), .ZN(n12165) );
  NAND2_X2 U11369 ( .A1(n12786), .A2(n12787), .ZN(n12169) );
  NAND2_X2 U11370 ( .A1(n11435), .A2(n11436), .ZN(n11643) );
  NAND2_X2 U11371 ( .A1(n12812), .A2(n12787), .ZN(n12199) );
  OAI21_X2 U11372 ( .B1(n25400), .B2(n26290), .A(n16353), .ZN(n16352) );
  OAI21_X2 U11373 ( .B1(n13032), .B2(n26293), .A(n16344), .ZN(n16343) );
  OAI21_X2 U11374 ( .B1(n15513), .B2(n15530), .A(n15536), .ZN(n15535) );
  NAND2_X2 U11375 ( .A1(n12812), .A2(n12789), .ZN(n12218) );
  NOR2_X2 U11376 ( .A1(n11788), .A2(n26303), .ZN(n11638) );
  NAND2_X2 U11377 ( .A1(n12788), .A2(n12789), .ZN(n12167) );
  INV_X4 U11378 ( .A(n12970), .ZN(n26509) );
  NAND2_X2 U11379 ( .A1(n11874), .A2(n24894), .ZN(n11801) );
  INV_X4 U11380 ( .A(n16210), .ZN(n26510) );
  AOI21_X2 U11381 ( .B1(n13078), .B2(n11634), .A(n26295), .ZN(n13076) );
  AOI21_X2 U11382 ( .B1(n25959), .B2(n11433), .A(n11435), .ZN(n11434) );
  OAI21_X2 U11383 ( .B1(n25253), .B2(n26293), .A(n13076), .ZN(n11400) );
  INV_X4 U11384 ( .A(n11813), .ZN(n26345) );
  INV_X4 U11385 ( .A(n11803), .ZN(n26342) );
  INV_X4 U11386 ( .A(n11806), .ZN(n26348) );
  INV_X4 U11387 ( .A(n10081), .ZN(n26130) );
  INV_X4 U11388 ( .A(n11809), .ZN(n26347) );
  AOI21_X2 U11389 ( .B1(n13069), .B2(n25956), .A(n26137), .ZN(n13068) );
  AOI22_X2 U11390 ( .A1(U7_DATA2_4), .A2(n26302), .B1(n26301), .B2(
        add_283_A_4_), .ZN(n13050) );
  AOI22_X2 U11391 ( .A1(U7_DATA2_3), .A2(n26302), .B1(n26301), .B2(
        add_283_A_3_), .ZN(n13051) );
  AOI22_X2 U11392 ( .A1(U7_DATA2_2), .A2(n26302), .B1(n26301), .B2(
        add_283_A_2_), .ZN(n13052) );
  AOI22_X2 U11393 ( .A1(U7_DATA2_1), .A2(n26302), .B1(n26301), .B2(
        add_283_A_1_), .ZN(n13053) );
  INV_X4 U11394 ( .A(n4890), .ZN(n25982) );
  INV_X4 U11395 ( .A(bvm__dut__data[3]), .ZN(n26131) );
  INV_X4 U11396 ( .A(bvm__dut__data[2]), .ZN(n26132) );
  INV_X4 U11397 ( .A(bvm__dut__data[1]), .ZN(n26133) );
  INV_X4 U11398 ( .A(bvm__dut__data[0]), .ZN(n26134) );
  OAI222_X2 U11399 ( .A1(n25901), .A2(n27403), .B1(n25899), .B2(n27467), .C1(
        n16811), .C2(n25898), .ZN(n15067) );
  OAI222_X2 U11400 ( .A1(n25902), .A2(n27404), .B1(n25900), .B2(n27468), .C1(
        n16774), .C2(n25898), .ZN(n15104) );
  OAI222_X2 U11401 ( .A1(n25901), .A2(n27402), .B1(n25900), .B2(n27466), .C1(
        n16848), .C2(n25897), .ZN(n15030) );
  OAI222_X2 U11402 ( .A1(n25901), .A2(n27400), .B1(n25899), .B2(n27464), .C1(
        n16922), .C2(n25898), .ZN(n14956) );
  OAI222_X2 U11403 ( .A1(n25902), .A2(n27401), .B1(n25899), .B2(n27465), .C1(
        n16885), .C2(n25897), .ZN(n14993) );
  OAI222_X2 U11404 ( .A1(n25901), .A2(n27399), .B1(n25900), .B2(n27463), .C1(
        n16959), .C2(n25897), .ZN(n14919) );
  OAI222_X2 U11405 ( .A1(n25902), .A2(n27362), .B1(n25900), .B2(n27426), .C1(
        n17144), .C2(n25898), .ZN(n14734) );
  OAI222_X2 U11406 ( .A1(n25902), .A2(n27361), .B1(n25900), .B2(n27425), .C1(
        n17181), .C2(n25898), .ZN(n14697) );
  OAI222_X2 U11407 ( .A1(n25902), .A2(n27360), .B1(n25900), .B2(n27424), .C1(
        n17218), .C2(n25898), .ZN(n14660) );
  OAI222_X2 U11408 ( .A1(n25902), .A2(n27359), .B1(n25900), .B2(n27423), .C1(
        n17255), .C2(n25898), .ZN(n14623) );
  OAI222_X2 U11409 ( .A1(n25902), .A2(n27358), .B1(n25900), .B2(n27422), .C1(
        n17292), .C2(n25898), .ZN(n14586) );
  OAI222_X2 U11410 ( .A1(n25902), .A2(n27357), .B1(n25900), .B2(n27421), .C1(
        n17329), .C2(n25898), .ZN(n14549) );
  OAI222_X2 U11411 ( .A1(n25902), .A2(n27356), .B1(n25900), .B2(n27420), .C1(
        n17366), .C2(n25898), .ZN(n14512) );
  OAI222_X2 U11412 ( .A1(n25902), .A2(n27355), .B1(n25899), .B2(n27419), .C1(
        n17403), .C2(n25898), .ZN(n14475) );
  OAI222_X2 U11413 ( .A1(n25901), .A2(n27354), .B1(n25900), .B2(n27418), .C1(
        n17440), .C2(n25897), .ZN(n14438) );
  OAI222_X2 U11414 ( .A1(n25901), .A2(n27353), .B1(n25899), .B2(n27417), .C1(
        n17477), .C2(n25897), .ZN(n14401) );
  OAI222_X2 U11415 ( .A1(n25901), .A2(n27352), .B1(n25900), .B2(n27416), .C1(
        n17514), .C2(n25897), .ZN(n14364) );
  OAI222_X2 U11416 ( .A1(n25901), .A2(n27351), .B1(n25899), .B2(n27415), .C1(
        n17551), .C2(n25897), .ZN(n14327) );
  OAI222_X2 U11417 ( .A1(n25901), .A2(n27378), .B1(n25900), .B2(n27442), .C1(
        n17736), .C2(n25897), .ZN(n14142) );
  OAI222_X2 U11418 ( .A1(n25901), .A2(n27377), .B1(n25899), .B2(n27441), .C1(
        n17773), .C2(n25897), .ZN(n14105) );
  OAI222_X2 U11419 ( .A1(n25901), .A2(n27376), .B1(n25900), .B2(n27440), .C1(
        n17810), .C2(n25897), .ZN(n14068) );
  OAI222_X2 U11420 ( .A1(n25901), .A2(n27375), .B1(n25900), .B2(n27439), .C1(
        n17847), .C2(n25897), .ZN(n14031) );
  OAI222_X2 U11421 ( .A1(n25901), .A2(n27374), .B1(n25900), .B2(n27438), .C1(
        n17884), .C2(n25897), .ZN(n13994) );
  OAI222_X2 U11422 ( .A1(n25902), .A2(n27373), .B1(n25900), .B2(n27437), .C1(
        n17921), .C2(n25897), .ZN(n13957) );
  OAI222_X2 U11423 ( .A1(n25901), .A2(n27372), .B1(n25900), .B2(n27436), .C1(
        n17958), .C2(n25897), .ZN(n13920) );
  OAI222_X2 U11424 ( .A1(n25901), .A2(n27371), .B1(n25900), .B2(n27435), .C1(
        n17995), .C2(n25898), .ZN(n13883) );
  OAI222_X2 U11425 ( .A1(n25902), .A2(n27370), .B1(n25900), .B2(n27434), .C1(
        n18032), .C2(n25897), .ZN(n13846) );
  OAI222_X2 U11426 ( .A1(n25902), .A2(n27369), .B1(n25900), .B2(n27433), .C1(
        n18069), .C2(n25897), .ZN(n13809) );
  OAI222_X2 U11427 ( .A1(n25901), .A2(n27368), .B1(n25900), .B2(n27432), .C1(
        n18106), .C2(n25897), .ZN(n13772) );
  OAI222_X2 U11428 ( .A1(n25902), .A2(n27367), .B1(n25900), .B2(n27431), .C1(
        n18143), .C2(n25897), .ZN(n13735) );
  OAI222_X2 U11429 ( .A1(n25901), .A2(n27394), .B1(n25899), .B2(n27458), .C1(
        n18328), .C2(n25897), .ZN(n13550) );
  OAI222_X2 U11430 ( .A1(n25901), .A2(n27393), .B1(n25899), .B2(n27457), .C1(
        n18365), .C2(n25898), .ZN(n13513) );
  OAI222_X2 U11431 ( .A1(n25902), .A2(n27392), .B1(n25899), .B2(n27456), .C1(
        n18402), .C2(n25897), .ZN(n13476) );
  OAI222_X2 U11432 ( .A1(n25902), .A2(n27391), .B1(n25899), .B2(n27455), .C1(
        n18439), .C2(n25897), .ZN(n13439) );
  OAI222_X2 U11433 ( .A1(n25901), .A2(n27390), .B1(n25899), .B2(n27454), .C1(
        n18476), .C2(n25898), .ZN(n13402) );
  OAI222_X2 U11434 ( .A1(n25901), .A2(n27389), .B1(n25899), .B2(n27453), .C1(
        n18513), .C2(n25897), .ZN(n13365) );
  OAI222_X2 U11435 ( .A1(n25902), .A2(n27388), .B1(n25899), .B2(n27452), .C1(
        n18550), .C2(n25897), .ZN(n13328) );
  OAI222_X2 U11436 ( .A1(n25902), .A2(n27387), .B1(n25899), .B2(n27451), .C1(
        n18587), .C2(n25898), .ZN(n13291) );
  OAI222_X2 U11437 ( .A1(n25901), .A2(n27386), .B1(n25899), .B2(n27450), .C1(
        n18624), .C2(n25898), .ZN(n13254) );
  OAI222_X2 U11438 ( .A1(n25901), .A2(n27385), .B1(n25899), .B2(n27449), .C1(
        n18661), .C2(n25897), .ZN(n13217) );
  OAI222_X2 U11439 ( .A1(n25902), .A2(n27384), .B1(n25899), .B2(n27448), .C1(
        n18698), .C2(n25897), .ZN(n13180) );
  OAI222_X2 U11440 ( .A1(n25902), .A2(n27383), .B1(n25899), .B2(n27447), .C1(
        n18735), .C2(n25898), .ZN(n13109) );
  INV_X4 U11441 ( .A(bvm__dut__data[6]), .ZN(n26277) );
  INV_X4 U11442 ( .A(bvm__dut__data[5]), .ZN(n26278) );
  INV_X4 U11443 ( .A(bvm__dut__data[4]), .ZN(n26279) );
  INV_X4 U11444 ( .A(bvm__dut__data[7]), .ZN(n26276) );
  INV_X4 U11445 ( .A(bvm__dut__data[8]), .ZN(n26275) );
  INV_X4 U11446 ( .A(bvm__dut__data[9]), .ZN(n26274) );
  INV_X4 U11447 ( .A(bvm__dut__data[10]), .ZN(n26273) );
  INV_X4 U11448 ( .A(bvm__dut__data[11]), .ZN(n26272) );
  INV_X4 U11449 ( .A(bvm__dut__data[12]), .ZN(n26271) );
  INV_X4 U11450 ( .A(bvm__dut__data[13]), .ZN(n26270) );
  INV_X4 U11451 ( .A(bvm__dut__data[14]), .ZN(n26269) );
  INV_X4 U11452 ( .A(bvm__dut__data[15]), .ZN(n26268) );
  NOR3_X2 U11453 ( .A1(n22427), .A2(n19349), .A3(n25958), .ZN(n11435) );
  OAI222_X2 U11454 ( .A1(n12180), .A2(n27879), .B1(n18795), .B2(n12182), .C1(
        n12183), .C2(n27959), .ZN(n12750) );
  OAI222_X2 U11455 ( .A1(n25884), .A2(n27595), .B1(n16785), .B2(n25881), .C1(
        n25880), .C2(n27787), .ZN(n15073) );
  OAI222_X2 U11456 ( .A1(n25883), .A2(n27596), .B1(n16748), .B2(n25882), .C1(
        n25879), .C2(n27788), .ZN(n15110) );
  OAI222_X2 U11457 ( .A1(n12180), .A2(n27884), .B1(n18980), .B2(n12182), .C1(
        n12183), .C2(n27964), .ZN(n12555) );
  OAI222_X2 U11458 ( .A1(n12180), .A2(n27880), .B1(n18832), .B2(n12182), .C1(
        n12183), .C2(n27960), .ZN(n12711) );
  OAI222_X2 U11459 ( .A1(n25883), .A2(n27594), .B1(n16822), .B2(n25881), .C1(
        n25879), .C2(n27786), .ZN(n15036) );
  OAI222_X2 U11460 ( .A1(n12180), .A2(n27881), .B1(n18869), .B2(n12182), .C1(
        n12183), .C2(n27961), .ZN(n12672) );
  OAI222_X2 U11461 ( .A1(n25884), .A2(n27592), .B1(n16896), .B2(n25882), .C1(
        n25880), .C2(n27784), .ZN(n14962) );
  OAI222_X2 U11462 ( .A1(n25883), .A2(n27593), .B1(n16859), .B2(n25881), .C1(
        n25880), .C2(n27785), .ZN(n14999) );
  OAI222_X2 U11463 ( .A1(n25884), .A2(n27591), .B1(n16933), .B2(n25881), .C1(
        n25879), .C2(n27783), .ZN(n14925) );
  OAI222_X2 U11464 ( .A1(n25884), .A2(n27554), .B1(n17118), .B2(n25882), .C1(
        n25880), .C2(n27746), .ZN(n14740) );
  OAI222_X2 U11465 ( .A1(n25883), .A2(n27553), .B1(n17155), .B2(n25882), .C1(
        n25880), .C2(n27745), .ZN(n14703) );
  OAI222_X2 U11466 ( .A1(n25884), .A2(n27552), .B1(n17192), .B2(n25882), .C1(
        n25879), .C2(n27744), .ZN(n14666) );
  OAI222_X2 U11467 ( .A1(n25884), .A2(n27551), .B1(n17229), .B2(n25882), .C1(
        n25879), .C2(n27743), .ZN(n14629) );
  OAI222_X2 U11468 ( .A1(n25883), .A2(n27550), .B1(n17266), .B2(n25882), .C1(
        n25880), .C2(n27742), .ZN(n14592) );
  OAI222_X2 U11469 ( .A1(n25883), .A2(n27549), .B1(n17303), .B2(n25882), .C1(
        n25879), .C2(n27741), .ZN(n14555) );
  OAI222_X2 U11470 ( .A1(n25884), .A2(n27548), .B1(n17340), .B2(n25882), .C1(
        n25880), .C2(n27740), .ZN(n14518) );
  OAI222_X2 U11471 ( .A1(n25883), .A2(n27547), .B1(n17377), .B2(n25882), .C1(
        n25879), .C2(n27739), .ZN(n14481) );
  OAI222_X2 U11472 ( .A1(n25883), .A2(n27546), .B1(n17414), .B2(n25882), .C1(
        n25879), .C2(n27738), .ZN(n14444) );
  OAI222_X2 U11473 ( .A1(n25884), .A2(n27545), .B1(n17451), .B2(n25881), .C1(
        n25880), .C2(n27737), .ZN(n14407) );
  OAI222_X2 U11474 ( .A1(n25883), .A2(n27544), .B1(n17488), .B2(n25881), .C1(
        n25879), .C2(n27736), .ZN(n14370) );
  OAI222_X2 U11475 ( .A1(n25884), .A2(n27543), .B1(n17525), .B2(n25881), .C1(
        n25880), .C2(n27735), .ZN(n14333) );
  OAI222_X2 U11476 ( .A1(n25884), .A2(n27570), .B1(n17710), .B2(n25882), .C1(
        n25879), .C2(n27762), .ZN(n14148) );
  OAI222_X2 U11477 ( .A1(n25883), .A2(n27569), .B1(n17747), .B2(n25881), .C1(
        n25880), .C2(n27761), .ZN(n14111) );
  OAI222_X2 U11478 ( .A1(n25884), .A2(n27568), .B1(n17784), .B2(n25881), .C1(
        n25879), .C2(n27760), .ZN(n14074) );
  OAI222_X2 U11479 ( .A1(n25883), .A2(n27567), .B1(n17821), .B2(n25881), .C1(
        n25880), .C2(n27759), .ZN(n14037) );
  OAI222_X2 U11480 ( .A1(n25884), .A2(n27566), .B1(n17858), .B2(n25881), .C1(
        n25880), .C2(n27758), .ZN(n14000) );
  OAI222_X2 U11481 ( .A1(n25884), .A2(n27565), .B1(n17895), .B2(n25881), .C1(
        n25880), .C2(n27757), .ZN(n13963) );
  OAI222_X2 U11482 ( .A1(n25884), .A2(n27564), .B1(n17932), .B2(n25881), .C1(
        n25880), .C2(n27756), .ZN(n13926) );
  OAI222_X2 U11483 ( .A1(n25884), .A2(n27563), .B1(n17969), .B2(n25881), .C1(
        n25880), .C2(n27755), .ZN(n13889) );
  OAI222_X2 U11484 ( .A1(n25884), .A2(n27562), .B1(n18006), .B2(n25881), .C1(
        n25880), .C2(n27754), .ZN(n13852) );
  OAI222_X2 U11485 ( .A1(n25884), .A2(n27561), .B1(n18043), .B2(n25881), .C1(
        n25880), .C2(n27753), .ZN(n13815) );
  OAI222_X2 U11486 ( .A1(n25884), .A2(n27560), .B1(n18080), .B2(n25881), .C1(
        n25880), .C2(n27752), .ZN(n13778) );
  OAI222_X2 U11487 ( .A1(n25884), .A2(n27559), .B1(n18117), .B2(n25881), .C1(
        n25880), .C2(n27751), .ZN(n13741) );
  OAI222_X2 U11488 ( .A1(n25883), .A2(n27586), .B1(n18302), .B2(n25882), .C1(
        n25879), .C2(n27778), .ZN(n13556) );
  OAI222_X2 U11489 ( .A1(n25883), .A2(n27585), .B1(n18339), .B2(n25882), .C1(
        n25879), .C2(n27777), .ZN(n13519) );
  OAI222_X2 U11490 ( .A1(n25883), .A2(n27584), .B1(n18376), .B2(n25881), .C1(
        n25879), .C2(n27776), .ZN(n13482) );
  OAI222_X2 U11491 ( .A1(n25883), .A2(n27583), .B1(n18413), .B2(n25881), .C1(
        n25879), .C2(n27775), .ZN(n13445) );
  OAI222_X2 U11492 ( .A1(n25883), .A2(n27582), .B1(n18450), .B2(n25882), .C1(
        n25879), .C2(n27774), .ZN(n13408) );
  OAI222_X2 U11493 ( .A1(n25883), .A2(n27581), .B1(n18487), .B2(n25882), .C1(
        n25879), .C2(n27773), .ZN(n13371) );
  OAI222_X2 U11494 ( .A1(n25883), .A2(n27580), .B1(n18524), .B2(n25881), .C1(
        n25879), .C2(n27772), .ZN(n13334) );
  OAI222_X2 U11495 ( .A1(n25883), .A2(n27579), .B1(n18561), .B2(n25881), .C1(
        n25879), .C2(n27771), .ZN(n13297) );
  OAI222_X2 U11496 ( .A1(n25883), .A2(n27578), .B1(n18598), .B2(n25882), .C1(
        n25879), .C2(n27770), .ZN(n13260) );
  OAI222_X2 U11497 ( .A1(n25883), .A2(n27577), .B1(n18635), .B2(n25882), .C1(
        n25879), .C2(n27769), .ZN(n13223) );
  OAI222_X2 U11498 ( .A1(n25883), .A2(n27576), .B1(n18672), .B2(n25881), .C1(
        n25879), .C2(n27768), .ZN(n13186) );
  OAI222_X2 U11499 ( .A1(n25883), .A2(n27575), .B1(n18709), .B2(n25881), .C1(
        n25879), .C2(n27767), .ZN(n13124) );
  OAI222_X2 U11500 ( .A1(n12180), .A2(n27878), .B1(n18758), .B2(n12182), .C1(
        n12183), .C2(n27958), .ZN(n12796) );
  OAI222_X2 U11501 ( .A1(n12180), .A2(n27882), .B1(n18906), .B2(n12182), .C1(
        n12183), .C2(n27962), .ZN(n12633) );
  OAI222_X2 U11502 ( .A1(n12180), .A2(n27883), .B1(n18943), .B2(n12182), .C1(
        n12183), .C2(n27963), .ZN(n12594) );
  OAI222_X2 U11503 ( .A1(n12180), .A2(n27885), .B1(n19017), .B2(n12182), .C1(
        n12183), .C2(n27965), .ZN(n12516) );
  OAI222_X2 U11504 ( .A1(n12180), .A2(n27886), .B1(n19054), .B2(n12182), .C1(
        n12183), .C2(n27966), .ZN(n12477) );
  OAI222_X2 U11505 ( .A1(n12180), .A2(n27887), .B1(n19091), .B2(n12182), .C1(
        n12183), .C2(n27967), .ZN(n12438) );
  OAI222_X2 U11506 ( .A1(n12180), .A2(n27888), .B1(n19128), .B2(n12182), .C1(
        n12183), .C2(n27968), .ZN(n12399) );
  OAI222_X2 U11507 ( .A1(n12180), .A2(n27889), .B1(n19165), .B2(n12182), .C1(
        n12183), .C2(n27969), .ZN(n12360) );
  OAI222_X2 U11508 ( .A1(n25901), .A2(n27406), .B1(n25900), .B2(n27470), .C1(
        n16700), .C2(n25897), .ZN(n15178) );
  OAI222_X2 U11509 ( .A1(n25884), .A2(n27598), .B1(n16674), .B2(n25882), .C1(
        n25879), .C2(n27790), .ZN(n15184) );
  OAI222_X2 U11510 ( .A1(n25901), .A2(n27410), .B1(n25899), .B2(n27474), .C1(
        n16552), .C2(n25897), .ZN(n15326) );
  OAI222_X2 U11511 ( .A1(n25901), .A2(n27409), .B1(n25899), .B2(n27473), .C1(
        n16589), .C2(n25898), .ZN(n15289) );
  OAI222_X2 U11512 ( .A1(n25902), .A2(n27408), .B1(n25899), .B2(n27472), .C1(
        n16626), .C2(n25897), .ZN(n15252) );
  OAI222_X2 U11513 ( .A1(n25902), .A2(n27407), .B1(n25900), .B2(n27471), .C1(
        n16663), .C2(n25898), .ZN(n15215) );
  OAI222_X2 U11514 ( .A1(n25902), .A2(n27405), .B1(n25899), .B2(n27469), .C1(
        n16737), .C2(n25898), .ZN(n15141) );
  OAI222_X2 U11515 ( .A1(n25902), .A2(n27366), .B1(n25900), .B2(n27430), .C1(
        n16996), .C2(n25898), .ZN(n14882) );
  OAI222_X2 U11516 ( .A1(n25902), .A2(n27365), .B1(n25900), .B2(n27429), .C1(
        n17033), .C2(n25898), .ZN(n14845) );
  OAI222_X2 U11517 ( .A1(n25902), .A2(n27364), .B1(n25899), .B2(n27428), .C1(
        n17070), .C2(n25898), .ZN(n14808) );
  OAI222_X2 U11518 ( .A1(n25902), .A2(n27363), .B1(n25899), .B2(n27427), .C1(
        n17107), .C2(n25898), .ZN(n14771) );
  OAI222_X2 U11519 ( .A1(n25901), .A2(n27382), .B1(n25900), .B2(n27446), .C1(
        n17588), .C2(n25897), .ZN(n14290) );
  OAI222_X2 U11520 ( .A1(n25901), .A2(n27381), .B1(n25899), .B2(n27445), .C1(
        n17625), .C2(n25897), .ZN(n14253) );
  OAI222_X2 U11521 ( .A1(n25901), .A2(n27380), .B1(n25899), .B2(n27444), .C1(
        n17662), .C2(n25897), .ZN(n14216) );
  OAI222_X2 U11522 ( .A1(n25901), .A2(n27379), .B1(n25900), .B2(n27443), .C1(
        n17699), .C2(n25897), .ZN(n14179) );
  OAI222_X2 U11523 ( .A1(n25901), .A2(n27398), .B1(n25900), .B2(n27462), .C1(
        n18180), .C2(n25897), .ZN(n13698) );
  OAI222_X2 U11524 ( .A1(n25902), .A2(n27397), .B1(n25900), .B2(n27461), .C1(
        n18217), .C2(n25897), .ZN(n13661) );
  OAI222_X2 U11525 ( .A1(n25901), .A2(n27396), .B1(n25900), .B2(n27460), .C1(
        n18254), .C2(n25897), .ZN(n13624) );
  OAI222_X2 U11526 ( .A1(n25901), .A2(n27395), .B1(n25899), .B2(n27459), .C1(
        n18291), .C2(n25898), .ZN(n13587) );
  OAI222_X2 U11527 ( .A1(n19217), .A2(n12215), .B1(n12216), .B2(n27938), .C1(
        n19216), .C2(n12218), .ZN(n12338) );
  OAI222_X2 U11528 ( .A1(n19254), .A2(n12215), .B1(n12216), .B2(n27939), .C1(
        n19253), .C2(n12218), .ZN(n12299) );
  OAI222_X2 U11529 ( .A1(n19291), .A2(n12215), .B1(n12216), .B2(n27940), .C1(
        n19290), .C2(n12218), .ZN(n12260) );
  OAI222_X2 U11530 ( .A1(n19328), .A2(n12215), .B1(n12216), .B2(n27941), .C1(
        n19327), .C2(n12218), .ZN(n12214) );
  AOI21_X2 U11531 ( .B1(n16185), .B2(n26501), .A(n22381), .ZN(n11487) );
  OAI222_X2 U11532 ( .A1(n18750), .A2(n11437), .B1(n12975), .B2(n12966), .C1(
        n22408), .C2(n25958), .ZN(n23269) );
  OAI222_X2 U11533 ( .A1(n18751), .A2(n11437), .B1(n12974), .B2(n12966), .C1(
        n22409), .C2(n25958), .ZN(n23268) );
  OAI222_X2 U11534 ( .A1(n18752), .A2(n11437), .B1(n26504), .B2(n12966), .C1(
        n22410), .C2(n25958), .ZN(n23267) );
  OAI222_X2 U11535 ( .A1(n18753), .A2(n11437), .B1(n12969), .B2(n12966), .C1(
        n22411), .C2(n25958), .ZN(n23266) );
  OAI222_X2 U11536 ( .A1(n18754), .A2(n11437), .B1(n12968), .B2(n12966), .C1(
        n22412), .C2(n25958), .ZN(n23265) );
  OAI222_X2 U11537 ( .A1(n18755), .A2(n11437), .B1(n12965), .B2(n12966), .C1(
        n22413), .C2(n25958), .ZN(n23264) );
  OAI222_X2 U11538 ( .A1(n15514), .A2(n15530), .B1(n12817), .B2(n15531), .C1(
        n22395), .C2(n26286), .ZN(n23516) );
  OAI222_X2 U11539 ( .A1(n12971), .A2(n16348), .B1(n16298), .B2(n26290), .C1(
        n22383), .C2(n26289), .ZN(n24814) );
  OAI222_X2 U11540 ( .A1(n22397), .A2(n15536), .B1(n15518), .B2(n15531), .C1(
        n15517), .C2(n15530), .ZN(n23518) );
  OAI222_X2 U11541 ( .A1(n26293), .A2(n26514), .B1(n16192), .B2(n16342), .C1(
        n22389), .C2(n16344), .ZN(n24812) );
  NOR4_X2 U11542 ( .A1(add_180_A_2_), .A2(add_180_A_1_), .A3(add_180_A_0_), 
        .A4(n22391), .ZN(n12813) );
  NAND4_X2 U11543 ( .A1(n11435), .A2(n22424), .A3(n24891), .A4(n25248), .ZN(
        n11649) );
  NOR4_X2 U11544 ( .A1(add_180_A_3_), .A2(add_180_A_1_), .A3(add_180_A_0_), 
        .A4(n22392), .ZN(n12812) );
  NAND4_X2 U11545 ( .A1(n11435), .A2(n22423), .A3(n24868), .A4(n25248), .ZN(
        n11651) );
  AOI22_X2 U11546 ( .A1(n11497), .A2(n16177), .B1(n11498), .B2(n26511), .ZN(
        n16180) );
  AOI21_X2 U11547 ( .B1(n16201), .B2(n11492), .A(n16202), .ZN(n16199) );
  NOR2_X2 U11548 ( .A1(add_283_A_2_), .A2(n22416), .ZN(n11196) );
  OAI222_X2 U11549 ( .A1(n18810), .A2(n12215), .B1(n12216), .B2(n27927), .C1(
        n18809), .C2(n12218), .ZN(n12767) );
  OAI222_X2 U11550 ( .A1(n18995), .A2(n12215), .B1(n12216), .B2(n27932), .C1(
        n18994), .C2(n12218), .ZN(n12572) );
  OAI222_X2 U11551 ( .A1(n18847), .A2(n12215), .B1(n12216), .B2(n27928), .C1(
        n18846), .C2(n12218), .ZN(n12728) );
  OAI222_X2 U11552 ( .A1(n18884), .A2(n12215), .B1(n12216), .B2(n27929), .C1(
        n18883), .C2(n12218), .ZN(n12689) );
  OAI222_X2 U11553 ( .A1(n17798), .A2(n25847), .B1(n17807), .B2(n25845), .C1(
        n17789), .C2(n25844), .ZN(n14092) );
  OAI222_X2 U11554 ( .A1(n17835), .A2(n25847), .B1(n17844), .B2(n25846), .C1(
        n17826), .C2(n25844), .ZN(n14055) );
  OAI222_X2 U11555 ( .A1(n17872), .A2(n25847), .B1(n17881), .B2(n25846), .C1(
        n17863), .C2(n25844), .ZN(n14018) );
  OAI222_X2 U11556 ( .A1(n17909), .A2(n25848), .B1(n17918), .B2(n25846), .C1(
        n17900), .C2(n25844), .ZN(n13981) );
  OAI222_X2 U11557 ( .A1(n17946), .A2(n25848), .B1(n17955), .B2(n25846), .C1(
        n17937), .C2(n25844), .ZN(n13944) );
  OAI222_X2 U11558 ( .A1(n17983), .A2(n25847), .B1(n17992), .B2(n25846), .C1(
        n17974), .C2(n25844), .ZN(n13907) );
  OAI222_X2 U11559 ( .A1(n18020), .A2(n25848), .B1(n18029), .B2(n25846), .C1(
        n18011), .C2(n25844), .ZN(n13870) );
  OAI222_X2 U11560 ( .A1(n18057), .A2(n25847), .B1(n18066), .B2(n25846), .C1(
        n18048), .C2(n25844), .ZN(n13833) );
  OAI222_X2 U11561 ( .A1(n18094), .A2(n25847), .B1(n18103), .B2(n25846), .C1(
        n18085), .C2(n25844), .ZN(n13796) );
  OAI222_X2 U11562 ( .A1(n18131), .A2(n25848), .B1(n18140), .B2(n25846), .C1(
        n18122), .C2(n25844), .ZN(n13759) );
  OAI222_X2 U11563 ( .A1(n18316), .A2(n25848), .B1(n18325), .B2(n25845), .C1(
        n18307), .C2(n25843), .ZN(n13574) );
  OAI222_X2 U11564 ( .A1(n18353), .A2(n25848), .B1(n18362), .B2(n25845), .C1(
        n18344), .C2(n25843), .ZN(n13537) );
  OAI222_X2 U11565 ( .A1(n18390), .A2(n25848), .B1(n18399), .B2(n25845), .C1(
        n18381), .C2(n25843), .ZN(n13500) );
  OAI222_X2 U11566 ( .A1(n18427), .A2(n25847), .B1(n18436), .B2(n25845), .C1(
        n18418), .C2(n25843), .ZN(n13463) );
  OAI222_X2 U11567 ( .A1(n18464), .A2(n25848), .B1(n18473), .B2(n25845), .C1(
        n18455), .C2(n25843), .ZN(n13426) );
  OAI222_X2 U11568 ( .A1(n18501), .A2(n25848), .B1(n18510), .B2(n25845), .C1(
        n18492), .C2(n25843), .ZN(n13389) );
  OAI222_X2 U11569 ( .A1(n18538), .A2(n25847), .B1(n18547), .B2(n25845), .C1(
        n18529), .C2(n25843), .ZN(n13352) );
  OAI222_X2 U11570 ( .A1(n18575), .A2(n25848), .B1(n18584), .B2(n25845), .C1(
        n18566), .C2(n25843), .ZN(n13315) );
  OAI222_X2 U11571 ( .A1(n18612), .A2(n25847), .B1(n18621), .B2(n25845), .C1(
        n18603), .C2(n25843), .ZN(n13278) );
  OAI222_X2 U11572 ( .A1(n18649), .A2(n25848), .B1(n18658), .B2(n25845), .C1(
        n18640), .C2(n25843), .ZN(n13241) );
  OAI222_X2 U11573 ( .A1(n18686), .A2(n25847), .B1(n18695), .B2(n25845), .C1(
        n18677), .C2(n25843), .ZN(n13204) );
  OAI222_X2 U11574 ( .A1(n18723), .A2(n25848), .B1(n18732), .B2(n25845), .C1(
        n18714), .C2(n25843), .ZN(n13160) );
  OAI222_X2 U11575 ( .A1(n18773), .A2(n12215), .B1(n12216), .B2(n27926), .C1(
        n18772), .C2(n12218), .ZN(n12823) );
  OAI222_X2 U11576 ( .A1(n18921), .A2(n12215), .B1(n12216), .B2(n27930), .C1(
        n18920), .C2(n12218), .ZN(n12650) );
  OAI222_X2 U11577 ( .A1(n18958), .A2(n12215), .B1(n12216), .B2(n27931), .C1(
        n18957), .C2(n12218), .ZN(n12611) );
  OAI222_X2 U11578 ( .A1(n19032), .A2(n12215), .B1(n12216), .B2(n27933), .C1(
        n19031), .C2(n12218), .ZN(n12533) );
  OAI222_X2 U11579 ( .A1(n19069), .A2(n12215), .B1(n12216), .B2(n27934), .C1(
        n19068), .C2(n12218), .ZN(n12494) );
  OAI222_X2 U11580 ( .A1(n19106), .A2(n12215), .B1(n12216), .B2(n27935), .C1(
        n19105), .C2(n12218), .ZN(n12455) );
  OAI222_X2 U11581 ( .A1(n19143), .A2(n12215), .B1(n12216), .B2(n27936), .C1(
        n19142), .C2(n12218), .ZN(n12416) );
  OAI222_X2 U11582 ( .A1(n19180), .A2(n12215), .B1(n12216), .B2(n27937), .C1(
        n19179), .C2(n12218), .ZN(n12377) );
  OAI222_X2 U11583 ( .A1(n25884), .A2(n27590), .B1(n18154), .B2(n25881), .C1(
        n25880), .C2(n27782), .ZN(n13704) );
  OAI222_X2 U11584 ( .A1(n18168), .A2(n25848), .B1(n18177), .B2(n25846), .C1(
        n18159), .C2(n25844), .ZN(n13722) );
  OAI222_X2 U11585 ( .A1(n25884), .A2(n27589), .B1(n18191), .B2(n25881), .C1(
        n25880), .C2(n27781), .ZN(n13667) );
  OAI222_X2 U11586 ( .A1(n18205), .A2(n25847), .B1(n18214), .B2(n25846), .C1(
        n18196), .C2(n25844), .ZN(n13685) );
  OAI222_X2 U11587 ( .A1(n25884), .A2(n27588), .B1(n18228), .B2(n25881), .C1(
        n25880), .C2(n27780), .ZN(n13630) );
  OAI222_X2 U11588 ( .A1(n18242), .A2(n25847), .B1(n18251), .B2(n25846), .C1(
        n18233), .C2(n25844), .ZN(n13648) );
  OAI222_X2 U11589 ( .A1(n25884), .A2(n27587), .B1(n18265), .B2(n25881), .C1(
        n25880), .C2(n27779), .ZN(n13593) );
  OAI222_X2 U11590 ( .A1(n18279), .A2(n25847), .B1(n18288), .B2(n25846), .C1(
        n18270), .C2(n25844), .ZN(n13611) );
  OAI222_X2 U11591 ( .A1(n16799), .A2(n25848), .B1(n16808), .B2(n25845), .C1(
        n16790), .C2(n25844), .ZN(n15091) );
  OAI222_X2 U11592 ( .A1(n16762), .A2(n25848), .B1(n16771), .B2(n25846), .C1(
        n16753), .C2(n25844), .ZN(n15128) );
  OAI222_X2 U11593 ( .A1(n16836), .A2(n25848), .B1(n16845), .B2(n25846), .C1(
        n16827), .C2(n25843), .ZN(n15054) );
  OAI222_X2 U11594 ( .A1(n16910), .A2(n25848), .B1(n16919), .B2(n25845), .C1(
        n16901), .C2(n25843), .ZN(n14980) );
  OAI222_X2 U11595 ( .A1(n16873), .A2(n25848), .B1(n16882), .B2(n25845), .C1(
        n16864), .C2(n25844), .ZN(n15017) );
  OAI222_X2 U11596 ( .A1(n16947), .A2(n25848), .B1(n16956), .B2(n25846), .C1(
        n16938), .C2(n25843), .ZN(n14943) );
  OAI222_X2 U11597 ( .A1(n17132), .A2(n25847), .B1(n17141), .B2(n25846), .C1(
        n17123), .C2(n25843), .ZN(n14758) );
  OAI222_X2 U11598 ( .A1(n17169), .A2(n25847), .B1(n17178), .B2(n25846), .C1(
        n17160), .C2(n25844), .ZN(n14721) );
  OAI222_X2 U11599 ( .A1(n17206), .A2(n25848), .B1(n17215), .B2(n25845), .C1(
        n17197), .C2(n25844), .ZN(n14684) );
  OAI222_X2 U11600 ( .A1(n17243), .A2(n25847), .B1(n17252), .B2(n25845), .C1(
        n17234), .C2(n25844), .ZN(n14647) );
  OAI222_X2 U11601 ( .A1(n17280), .A2(n25848), .B1(n17289), .B2(n25846), .C1(
        n17271), .C2(n25843), .ZN(n14610) );
  OAI222_X2 U11602 ( .A1(n17317), .A2(n25847), .B1(n17326), .B2(n25845), .C1(
        n17308), .C2(n25844), .ZN(n14573) );
  OAI222_X2 U11603 ( .A1(n17354), .A2(n25847), .B1(n17363), .B2(n25846), .C1(
        n17345), .C2(n25843), .ZN(n14536) );
  OAI222_X2 U11604 ( .A1(n17391), .A2(n25847), .B1(n17400), .B2(n25845), .C1(
        n17382), .C2(n25844), .ZN(n14499) );
  OAI222_X2 U11605 ( .A1(n17428), .A2(n25847), .B1(n17437), .B2(n25845), .C1(
        n17419), .C2(n25844), .ZN(n14462) );
  OAI222_X2 U11606 ( .A1(n17465), .A2(n25847), .B1(n17474), .B2(n25846), .C1(
        n17456), .C2(n25843), .ZN(n14425) );
  OAI222_X2 U11607 ( .A1(n17502), .A2(n25847), .B1(n17511), .B2(n25845), .C1(
        n17493), .C2(n25844), .ZN(n14388) );
  OAI222_X2 U11608 ( .A1(n17539), .A2(n25847), .B1(n17548), .B2(n25846), .C1(
        n17530), .C2(n25843), .ZN(n14351) );
  OAI222_X2 U11609 ( .A1(n17724), .A2(n25847), .B1(n17733), .B2(n25845), .C1(
        n17715), .C2(n25844), .ZN(n14166) );
  OAI222_X2 U11610 ( .A1(n17761), .A2(n25847), .B1(n17770), .B2(n25846), .C1(
        n17752), .C2(n25844), .ZN(n14129) );
  OAI222_X2 U11611 ( .A1(n16688), .A2(n25848), .B1(n16697), .B2(n25846), .C1(
        n16679), .C2(n25844), .ZN(n15202) );
  OAI222_X2 U11612 ( .A1(n25884), .A2(n27606), .B1(n16378), .B2(n25882), .C1(
        n25879), .C2(n27798), .ZN(n15485) );
  OAI222_X2 U11613 ( .A1(n16392), .A2(n25847), .B1(n16401), .B2(n25846), .C1(
        n16383), .C2(n25843), .ZN(n15504) );
  OAI222_X2 U11614 ( .A1(n25884), .A2(n27605), .B1(n16415), .B2(n25882), .C1(
        n25879), .C2(n27797), .ZN(n15443) );
  OAI222_X2 U11615 ( .A1(n16429), .A2(n25847), .B1(n16438), .B2(n25845), .C1(
        n16420), .C2(n25843), .ZN(n15461) );
  OAI222_X2 U11616 ( .A1(n25883), .A2(n27604), .B1(n16452), .B2(n25882), .C1(
        n25880), .C2(n27796), .ZN(n15406) );
  OAI222_X2 U11617 ( .A1(n16466), .A2(n25848), .B1(n16475), .B2(n25845), .C1(
        n16457), .C2(n25843), .ZN(n15424) );
  OAI222_X2 U11618 ( .A1(n25883), .A2(n27603), .B1(n16489), .B2(n25882), .C1(
        n25880), .C2(n27795), .ZN(n15369) );
  OAI222_X2 U11619 ( .A1(n16503), .A2(n25848), .B1(n16512), .B2(n25846), .C1(
        n16494), .C2(n25844), .ZN(n15387) );
  OAI222_X2 U11620 ( .A1(n25884), .A2(n27602), .B1(n16526), .B2(n25881), .C1(
        n25880), .C2(n27794), .ZN(n15332) );
  OAI222_X2 U11621 ( .A1(n16540), .A2(n25848), .B1(n16549), .B2(n25845), .C1(
        n16531), .C2(n25844), .ZN(n15350) );
  OAI222_X2 U11622 ( .A1(n25883), .A2(n27601), .B1(n16563), .B2(n25882), .C1(
        n25879), .C2(n27793), .ZN(n15295) );
  OAI222_X2 U11623 ( .A1(n16577), .A2(n25848), .B1(n16586), .B2(n25846), .C1(
        n16568), .C2(n25843), .ZN(n15313) );
  OAI222_X2 U11624 ( .A1(n25883), .A2(n27600), .B1(n16600), .B2(n25881), .C1(
        n25880), .C2(n27792), .ZN(n15258) );
  OAI222_X2 U11625 ( .A1(n16614), .A2(n25848), .B1(n16623), .B2(n25846), .C1(
        n16605), .C2(n25844), .ZN(n15276) );
  OAI222_X2 U11626 ( .A1(n25884), .A2(n27599), .B1(n16637), .B2(n25881), .C1(
        n25879), .C2(n27791), .ZN(n15221) );
  OAI222_X2 U11627 ( .A1(n16651), .A2(n25848), .B1(n16660), .B2(n25845), .C1(
        n16642), .C2(n25843), .ZN(n15239) );
  OAI222_X2 U11628 ( .A1(n25883), .A2(n27597), .B1(n16711), .B2(n25881), .C1(
        n25880), .C2(n27789), .ZN(n15147) );
  OAI222_X2 U11629 ( .A1(n16725), .A2(n25848), .B1(n16734), .B2(n25845), .C1(
        n16716), .C2(n25844), .ZN(n15165) );
  OAI222_X2 U11630 ( .A1(n25884), .A2(n27558), .B1(n16970), .B2(n25882), .C1(
        n25879), .C2(n27750), .ZN(n14888) );
  OAI222_X2 U11631 ( .A1(n16984), .A2(n25848), .B1(n16993), .B2(n25846), .C1(
        n16975), .C2(n25843), .ZN(n14906) );
  OAI222_X2 U11632 ( .A1(n25883), .A2(n27557), .B1(n17007), .B2(n25882), .C1(
        n25880), .C2(n27749), .ZN(n14851) );
  OAI222_X2 U11633 ( .A1(n17021), .A2(n25847), .B1(n17030), .B2(n25845), .C1(
        n17012), .C2(n25844), .ZN(n14869) );
  OAI222_X2 U11634 ( .A1(n25883), .A2(n27556), .B1(n17044), .B2(n25882), .C1(
        n25879), .C2(n27748), .ZN(n14814) );
  OAI222_X2 U11635 ( .A1(n17058), .A2(n25847), .B1(n17067), .B2(n25846), .C1(
        n17049), .C2(n25844), .ZN(n14832) );
  OAI222_X2 U11636 ( .A1(n25884), .A2(n27555), .B1(n17081), .B2(n25882), .C1(
        n25880), .C2(n27747), .ZN(n14777) );
  OAI222_X2 U11637 ( .A1(n17095), .A2(n25848), .B1(n17104), .B2(n25845), .C1(
        n17086), .C2(n25844), .ZN(n14795) );
  OAI222_X2 U11638 ( .A1(n25883), .A2(n27574), .B1(n17562), .B2(n25882), .C1(
        n25879), .C2(n27766), .ZN(n14296) );
  OAI222_X2 U11639 ( .A1(n17576), .A2(n25847), .B1(n17585), .B2(n25845), .C1(
        n17567), .C2(n25843), .ZN(n14314) );
  OAI222_X2 U11640 ( .A1(n25884), .A2(n27573), .B1(n17599), .B2(n25882), .C1(
        n25880), .C2(n27765), .ZN(n14259) );
  OAI222_X2 U11641 ( .A1(n17613), .A2(n25847), .B1(n17622), .B2(n25846), .C1(
        n17604), .C2(n25844), .ZN(n14277) );
  OAI222_X2 U11642 ( .A1(n25884), .A2(n27572), .B1(n17636), .B2(n25881), .C1(
        n25880), .C2(n27764), .ZN(n14222) );
  OAI222_X2 U11643 ( .A1(n17650), .A2(n25847), .B1(n17659), .B2(n25845), .C1(
        n17641), .C2(n25843), .ZN(n14240) );
  OAI222_X2 U11644 ( .A1(n25883), .A2(n27571), .B1(n17673), .B2(n25881), .C1(
        n25879), .C2(n27763), .ZN(n14185) );
  OAI222_X2 U11645 ( .A1(n17687), .A2(n25847), .B1(n17696), .B2(n25846), .C1(
        n17678), .C2(n25843), .ZN(n14203) );
  OAI222_X2 U11646 ( .A1(n12180), .A2(n27890), .B1(n19202), .B2(n12182), .C1(
        n12183), .C2(n27970), .ZN(n12321) );
  OAI222_X2 U11647 ( .A1(n12180), .A2(n27891), .B1(n19239), .B2(n12182), .C1(
        n12183), .C2(n27971), .ZN(n12282) );
  OAI222_X2 U11648 ( .A1(n12180), .A2(n27892), .B1(n19276), .B2(n12182), .C1(
        n12183), .C2(n27972), .ZN(n12243) );
  OAI222_X2 U11649 ( .A1(n12180), .A2(n27893), .B1(n19313), .B2(n12182), .C1(
        n12183), .C2(n27973), .ZN(n12179) );
  OAI222_X2 U11650 ( .A1(n25866), .A2(n26992), .B1(n25864), .B2(n26800), .C1(
        n25861), .C2(n26928), .ZN(n14085) );
  OAI222_X2 U11651 ( .A1(n25865), .A2(n26991), .B1(n25864), .B2(n26799), .C1(
        n25862), .C2(n26927), .ZN(n14048) );
  OAI222_X2 U11652 ( .A1(n25866), .A2(n26990), .B1(n25864), .B2(n26798), .C1(
        n25862), .C2(n26926), .ZN(n14011) );
  OAI222_X2 U11653 ( .A1(n25866), .A2(n26989), .B1(n25864), .B2(n26797), .C1(
        n25862), .C2(n26925), .ZN(n13974) );
  OAI222_X2 U11654 ( .A1(n25866), .A2(n26988), .B1(n25864), .B2(n26796), .C1(
        n25862), .C2(n26924), .ZN(n13937) );
  OAI222_X2 U11655 ( .A1(n25866), .A2(n26987), .B1(n25864), .B2(n26795), .C1(
        n25862), .C2(n26923), .ZN(n13900) );
  OAI222_X2 U11656 ( .A1(n25866), .A2(n26986), .B1(n25864), .B2(n26794), .C1(
        n25862), .C2(n26922), .ZN(n13863) );
  OAI222_X2 U11657 ( .A1(n25866), .A2(n26985), .B1(n25864), .B2(n26793), .C1(
        n25862), .C2(n26921), .ZN(n13826) );
  OAI222_X2 U11658 ( .A1(n25866), .A2(n26984), .B1(n25864), .B2(n26792), .C1(
        n25862), .C2(n26920), .ZN(n13789) );
  OAI222_X2 U11659 ( .A1(n25866), .A2(n26983), .B1(n25864), .B2(n26791), .C1(
        n25862), .C2(n26919), .ZN(n13752) );
  OAI222_X2 U11660 ( .A1(n25865), .A2(n27010), .B1(n25863), .B2(n26818), .C1(
        n25861), .C2(n26946), .ZN(n13567) );
  OAI222_X2 U11661 ( .A1(n25865), .A2(n27009), .B1(n25863), .B2(n26817), .C1(
        n25861), .C2(n26945), .ZN(n13530) );
  OAI222_X2 U11662 ( .A1(n25865), .A2(n27008), .B1(n25863), .B2(n26816), .C1(
        n25861), .C2(n26944), .ZN(n13493) );
  OAI222_X2 U11663 ( .A1(n25865), .A2(n27007), .B1(n25863), .B2(n26815), .C1(
        n25861), .C2(n26943), .ZN(n13456) );
  OAI222_X2 U11664 ( .A1(n25865), .A2(n27006), .B1(n25863), .B2(n26814), .C1(
        n25861), .C2(n26942), .ZN(n13419) );
  OAI222_X2 U11665 ( .A1(n25865), .A2(n27005), .B1(n25863), .B2(n26813), .C1(
        n25861), .C2(n26941), .ZN(n13382) );
  OAI222_X2 U11666 ( .A1(n25865), .A2(n27004), .B1(n25863), .B2(n26812), .C1(
        n25861), .C2(n26940), .ZN(n13345) );
  OAI222_X2 U11667 ( .A1(n25865), .A2(n27003), .B1(n25863), .B2(n26811), .C1(
        n25861), .C2(n26939), .ZN(n13308) );
  OAI222_X2 U11668 ( .A1(n25865), .A2(n27002), .B1(n25863), .B2(n26810), .C1(
        n25861), .C2(n26938), .ZN(n13271) );
  OAI222_X2 U11669 ( .A1(n25865), .A2(n27001), .B1(n25863), .B2(n26809), .C1(
        n25861), .C2(n26937), .ZN(n13234) );
  OAI222_X2 U11670 ( .A1(n25865), .A2(n27000), .B1(n25863), .B2(n26808), .C1(
        n25861), .C2(n26936), .ZN(n13197) );
  OAI222_X2 U11671 ( .A1(n25865), .A2(n26999), .B1(n25863), .B2(n26807), .C1(
        n25861), .C2(n26935), .ZN(n13144) );
  OAI222_X2 U11672 ( .A1(n25866), .A2(n27014), .B1(n25864), .B2(n26822), .C1(
        n25862), .C2(n26950), .ZN(n13715) );
  OAI222_X2 U11673 ( .A1(n25866), .A2(n27013), .B1(n25864), .B2(n26821), .C1(
        n25862), .C2(n26949), .ZN(n13678) );
  OAI222_X2 U11674 ( .A1(n25866), .A2(n27012), .B1(n25864), .B2(n26820), .C1(
        n25862), .C2(n26948), .ZN(n13641) );
  OAI222_X2 U11675 ( .A1(n25866), .A2(n27011), .B1(n25863), .B2(n26819), .C1(
        n25862), .C2(n26947), .ZN(n13604) );
  OAI222_X2 U11676 ( .A1(n25866), .A2(n27019), .B1(n25863), .B2(n26827), .C1(
        n25862), .C2(n26955), .ZN(n15084) );
  OAI222_X2 U11677 ( .A1(n25866), .A2(n27020), .B1(n25864), .B2(n26828), .C1(
        n25862), .C2(n26956), .ZN(n15121) );
  OAI222_X2 U11678 ( .A1(n25865), .A2(n27018), .B1(n25864), .B2(n26826), .C1(
        n25861), .C2(n26954), .ZN(n15047) );
  OAI222_X2 U11679 ( .A1(n25865), .A2(n27016), .B1(n25863), .B2(n26824), .C1(
        n25861), .C2(n26952), .ZN(n14973) );
  OAI222_X2 U11680 ( .A1(n25866), .A2(n27017), .B1(n25864), .B2(n26825), .C1(
        n25862), .C2(n26953), .ZN(n15010) );
  OAI222_X2 U11681 ( .A1(n25865), .A2(n27015), .B1(n25864), .B2(n26823), .C1(
        n25861), .C2(n26951), .ZN(n14936) );
  OAI222_X2 U11682 ( .A1(n25865), .A2(n26978), .B1(n25864), .B2(n26786), .C1(
        n25862), .C2(n26914), .ZN(n14751) );
  OAI222_X2 U11683 ( .A1(n25865), .A2(n26977), .B1(n25863), .B2(n26785), .C1(
        n25862), .C2(n26913), .ZN(n14714) );
  OAI222_X2 U11684 ( .A1(n25866), .A2(n26976), .B1(n25863), .B2(n26784), .C1(
        n25861), .C2(n26912), .ZN(n14677) );
  OAI222_X2 U11685 ( .A1(n25866), .A2(n26975), .B1(n25864), .B2(n26783), .C1(
        n25861), .C2(n26911), .ZN(n14640) );
  OAI222_X2 U11686 ( .A1(n25865), .A2(n26974), .B1(n25863), .B2(n26782), .C1(
        n25862), .C2(n26910), .ZN(n14603) );
  OAI222_X2 U11687 ( .A1(n25866), .A2(n26973), .B1(n25864), .B2(n26781), .C1(
        n25861), .C2(n26909), .ZN(n14566) );
  OAI222_X2 U11688 ( .A1(n25865), .A2(n26972), .B1(n25863), .B2(n26780), .C1(
        n25862), .C2(n26908), .ZN(n14529) );
  OAI222_X2 U11689 ( .A1(n25866), .A2(n26971), .B1(n25864), .B2(n26779), .C1(
        n25861), .C2(n26907), .ZN(n14492) );
  OAI222_X2 U11690 ( .A1(n25865), .A2(n26970), .B1(n25863), .B2(n26778), .C1(
        n25861), .C2(n26906), .ZN(n14455) );
  OAI222_X2 U11691 ( .A1(n25866), .A2(n26969), .B1(n25864), .B2(n26777), .C1(
        n25862), .C2(n26905), .ZN(n14418) );
  OAI222_X2 U11692 ( .A1(n25865), .A2(n26968), .B1(n25863), .B2(n26776), .C1(
        n25861), .C2(n26904), .ZN(n14381) );
  OAI222_X2 U11693 ( .A1(n25866), .A2(n26967), .B1(n25864), .B2(n26775), .C1(
        n25862), .C2(n26903), .ZN(n14344) );
  OAI222_X2 U11694 ( .A1(n25866), .A2(n26994), .B1(n25863), .B2(n26802), .C1(
        n25861), .C2(n26930), .ZN(n14159) );
  OAI222_X2 U11695 ( .A1(n25865), .A2(n26993), .B1(n25864), .B2(n26801), .C1(
        n25862), .C2(n26929), .ZN(n14122) );
  OAI222_X2 U11696 ( .A1(n25866), .A2(n27022), .B1(n25864), .B2(n26830), .C1(
        n25862), .C2(n26958), .ZN(n15195) );
  OAI222_X2 U11697 ( .A1(n25865), .A2(n27030), .B1(n25863), .B2(n26838), .C1(
        n25862), .C2(n26966), .ZN(n15497) );
  OAI222_X2 U11698 ( .A1(n25865), .A2(n27029), .B1(n25864), .B2(n26837), .C1(
        n25861), .C2(n26965), .ZN(n15454) );
  OAI222_X2 U11699 ( .A1(n25866), .A2(n27028), .B1(n25863), .B2(n26836), .C1(
        n25862), .C2(n26964), .ZN(n15417) );
  OAI222_X2 U11700 ( .A1(n25865), .A2(n27027), .B1(n25864), .B2(n26835), .C1(
        n25861), .C2(n26963), .ZN(n15380) );
  OAI222_X2 U11701 ( .A1(n25865), .A2(n27026), .B1(n25864), .B2(n26834), .C1(
        n25861), .C2(n26962), .ZN(n15343) );
  OAI222_X2 U11702 ( .A1(n25865), .A2(n27025), .B1(n25864), .B2(n26833), .C1(
        n25861), .C2(n26961), .ZN(n15306) );
  OAI222_X2 U11703 ( .A1(n25866), .A2(n27024), .B1(n25863), .B2(n26832), .C1(
        n25862), .C2(n26960), .ZN(n15269) );
  OAI222_X2 U11704 ( .A1(n25866), .A2(n27023), .B1(n25864), .B2(n26831), .C1(
        n25862), .C2(n26959), .ZN(n15232) );
  OAI222_X2 U11705 ( .A1(n25865), .A2(n27021), .B1(n25863), .B2(n26829), .C1(
        n25861), .C2(n26957), .ZN(n15158) );
  OAI222_X2 U11706 ( .A1(n25866), .A2(n26982), .B1(n25863), .B2(n26790), .C1(
        n25861), .C2(n26918), .ZN(n14899) );
  OAI222_X2 U11707 ( .A1(n25865), .A2(n26981), .B1(n25864), .B2(n26789), .C1(
        n25862), .C2(n26917), .ZN(n14862) );
  OAI222_X2 U11708 ( .A1(n25865), .A2(n26980), .B1(n25863), .B2(n26788), .C1(
        n25862), .C2(n26916), .ZN(n14825) );
  OAI222_X2 U11709 ( .A1(n25865), .A2(n26979), .B1(n25863), .B2(n26787), .C1(
        n25861), .C2(n26915), .ZN(n14788) );
  OAI222_X2 U11710 ( .A1(n25866), .A2(n26998), .B1(n25863), .B2(n26806), .C1(
        n25861), .C2(n26934), .ZN(n14307) );
  OAI222_X2 U11711 ( .A1(n25866), .A2(n26997), .B1(n25863), .B2(n26805), .C1(
        n25862), .C2(n26933), .ZN(n14270) );
  OAI222_X2 U11712 ( .A1(n25866), .A2(n26996), .B1(n25864), .B2(n26804), .C1(
        n25861), .C2(n26932), .ZN(n14233) );
  OAI222_X2 U11713 ( .A1(n25866), .A2(n26995), .B1(n25864), .B2(n26803), .C1(
        n25862), .C2(n26931), .ZN(n14196) );
  OAI222_X2 U11714 ( .A1(n18827), .A2(n12199), .B1(n18828), .B2(n12200), .C1(
        n12201), .C2(n27831), .ZN(n12760) );
  OAI222_X2 U11715 ( .A1(n19012), .A2(n12199), .B1(n19013), .B2(n12200), .C1(
        n12201), .C2(n27836), .ZN(n12565) );
  OAI222_X2 U11716 ( .A1(n18864), .A2(n12199), .B1(n18865), .B2(n12200), .C1(
        n12201), .C2(n27832), .ZN(n12721) );
  OAI222_X2 U11717 ( .A1(n18901), .A2(n12199), .B1(n18902), .B2(n12200), .C1(
        n12201), .C2(n27833), .ZN(n12682) );
  OAI222_X2 U11718 ( .A1(n12165), .A2(n28087), .B1(n12167), .B2(n28007), .C1(
        n18823), .C2(n12169), .ZN(n12744) );
  OAI222_X2 U11719 ( .A1(n12165), .A2(n28092), .B1(n12167), .B2(n28012), .C1(
        n19008), .C2(n12169), .ZN(n12549) );
  OAI222_X2 U11720 ( .A1(n12165), .A2(n28088), .B1(n12167), .B2(n28008), .C1(
        n18860), .C2(n12169), .ZN(n12705) );
  OAI222_X2 U11721 ( .A1(n12165), .A2(n28089), .B1(n12167), .B2(n28009), .C1(
        n18897), .C2(n12169), .ZN(n12666) );
  OAI222_X2 U11722 ( .A1(n18790), .A2(n12199), .B1(n18791), .B2(n12200), .C1(
        n12201), .C2(n27830), .ZN(n12808) );
  OAI222_X2 U11723 ( .A1(n18938), .A2(n12199), .B1(n18939), .B2(n12200), .C1(
        n12201), .C2(n27834), .ZN(n12643) );
  OAI222_X2 U11724 ( .A1(n18975), .A2(n12199), .B1(n18976), .B2(n12200), .C1(
        n12201), .C2(n27835), .ZN(n12604) );
  OAI222_X2 U11725 ( .A1(n19049), .A2(n12199), .B1(n19050), .B2(n12200), .C1(
        n12201), .C2(n27837), .ZN(n12526) );
  OAI222_X2 U11726 ( .A1(n19086), .A2(n12199), .B1(n19087), .B2(n12200), .C1(
        n12201), .C2(n27838), .ZN(n12487) );
  OAI222_X2 U11727 ( .A1(n19123), .A2(n12199), .B1(n19124), .B2(n12200), .C1(
        n12201), .C2(n27839), .ZN(n12448) );
  OAI222_X2 U11728 ( .A1(n19160), .A2(n12199), .B1(n19161), .B2(n12200), .C1(
        n12201), .C2(n27840), .ZN(n12409) );
  OAI222_X2 U11729 ( .A1(n19197), .A2(n12199), .B1(n19198), .B2(n12200), .C1(
        n12201), .C2(n27841), .ZN(n12370) );
  OAI222_X2 U11730 ( .A1(n12165), .A2(n28086), .B1(n12167), .B2(n28006), .C1(
        n18786), .C2(n12169), .ZN(n12783) );
  OAI222_X2 U11731 ( .A1(n12165), .A2(n28090), .B1(n12167), .B2(n28010), .C1(
        n18934), .C2(n12169), .ZN(n12627) );
  OAI222_X2 U11732 ( .A1(n12165), .A2(n28091), .B1(n12167), .B2(n28011), .C1(
        n18971), .C2(n12169), .ZN(n12588) );
  OAI222_X2 U11733 ( .A1(n12165), .A2(n28093), .B1(n12167), .B2(n28013), .C1(
        n19045), .C2(n12169), .ZN(n12510) );
  OAI222_X2 U11734 ( .A1(n12165), .A2(n28094), .B1(n12167), .B2(n28014), .C1(
        n19082), .C2(n12169), .ZN(n12471) );
  OAI222_X2 U11735 ( .A1(n12165), .A2(n28095), .B1(n12167), .B2(n28015), .C1(
        n19119), .C2(n12169), .ZN(n12432) );
  OAI222_X2 U11736 ( .A1(n12165), .A2(n28096), .B1(n12167), .B2(n28016), .C1(
        n19156), .C2(n12169), .ZN(n12393) );
  OAI222_X2 U11737 ( .A1(n12165), .A2(n28097), .B1(n12167), .B2(n28017), .C1(
        n19193), .C2(n12169), .ZN(n12354) );
  OAI222_X2 U11738 ( .A1(n19234), .A2(n12199), .B1(n19235), .B2(n12200), .C1(
        n12201), .C2(n27842), .ZN(n12331) );
  OAI222_X2 U11739 ( .A1(n19271), .A2(n12199), .B1(n19272), .B2(n12200), .C1(
        n12201), .C2(n27843), .ZN(n12292) );
  OAI222_X2 U11740 ( .A1(n19308), .A2(n12199), .B1(n19309), .B2(n12200), .C1(
        n12201), .C2(n27844), .ZN(n12253) );
  OAI222_X2 U11741 ( .A1(n19345), .A2(n12199), .B1(n19346), .B2(n12200), .C1(
        n12201), .C2(n27845), .ZN(n12198) );
  OAI222_X2 U11742 ( .A1(n25902), .A2(n27414), .B1(n25900), .B2(n27478), .C1(
        n16404), .C2(n25898), .ZN(n15474) );
  OAI222_X2 U11743 ( .A1(n25901), .A2(n27413), .B1(n25899), .B2(n27477), .C1(
        n16441), .C2(n25898), .ZN(n15437) );
  OAI222_X2 U11744 ( .A1(n25902), .A2(n27412), .B1(n25900), .B2(n27476), .C1(
        n16478), .C2(n25898), .ZN(n15400) );
  OAI222_X2 U11745 ( .A1(n25901), .A2(n27411), .B1(n25900), .B2(n27475), .C1(
        n16515), .C2(n25898), .ZN(n15363) );
  OAI222_X2 U11746 ( .A1(n12165), .A2(n28098), .B1(n12167), .B2(n28018), .C1(
        n19230), .C2(n12169), .ZN(n12315) );
  OAI222_X2 U11747 ( .A1(n12165), .A2(n28099), .B1(n12167), .B2(n28019), .C1(
        n19267), .C2(n12169), .ZN(n12276) );
  OAI222_X2 U11748 ( .A1(n12165), .A2(n28100), .B1(n12167), .B2(n28020), .C1(
        n19304), .C2(n12169), .ZN(n12237) );
  OAI222_X2 U11749 ( .A1(n12165), .A2(n28101), .B1(n12167), .B2(n28021), .C1(
        n19341), .C2(n12169), .ZN(n12164) );
  NOR2_X2 U11750 ( .A1(add_283_A_3_), .A2(n22417), .ZN(n11195) );
  OAI21_X2 U11751 ( .B1(n16207), .B2(n11491), .A(n26515), .ZN(n16211) );
  AOI22_X2 U11752 ( .A1(n16194), .A2(n11491), .B1(n22387), .B2(n26498), .ZN(
        n16193) );
  AOI21_X2 U11753 ( .B1(n11487), .B2(n16178), .A(n16179), .ZN(n16189) );
  AOI21_X2 U11754 ( .B1(n22423), .B2(n11634), .A(n16361), .ZN(n16360) );
  AOI21_X2 U11755 ( .B1(n11634), .B2(n22427), .A(n16346), .ZN(n16364) );
  OAI21_X2 U11756 ( .B1(n22399), .B2(n26350), .A(n11634), .ZN(n13075) );
  AOI21_X2 U11757 ( .B1(n22394), .B2(n15538), .A(n15537), .ZN(n15545) );
  AOI21_X2 U11758 ( .B1(n22386), .B2(n16347), .A(n16346), .ZN(n16353) );
  AOI21_X2 U11759 ( .B1(n22406), .B2(n13085), .A(n26295), .ZN(n13091) );
  AOI21_X2 U11760 ( .B1(n26507), .B2(n16196), .A(n12975), .ZN(n16200) );
  OAI211_X2 U11761 ( .C1(n16367), .C2(n11487), .A(n11488), .B(n11489), .ZN(
        n21419) );
  AOI21_X2 U11762 ( .B1(n15538), .B2(n22392), .A(n15541), .ZN(n15540) );
  OAI21_X2 U11763 ( .B1(n22392), .B2(n26284), .A(n15543), .ZN(n23521) );
  OAI21_X2 U11764 ( .B1(n22384), .B2(n26289), .A(n16351), .ZN(n24815) );
  OAI21_X2 U11765 ( .B1(n13060), .B2(n26296), .A(add_1445_B_9_), .ZN(n13057)
         );
  OAI21_X2 U11766 ( .B1(n16177), .B2(n16178), .A(n16179), .ZN(n16176) );
  OAI21_X2 U11767 ( .B1(n13081), .B2(n26136), .A(n13083), .ZN(n23447) );
  AOI21_X2 U11768 ( .B1(n13085), .B2(n22404), .A(n13086), .ZN(n13081) );
  OAI21_X2 U11769 ( .B1(n18746), .B2(n11437), .A(n11440), .ZN(n21154) );
  OAI21_X2 U11770 ( .B1(n18747), .B2(n11437), .A(n11439), .ZN(n21153) );
  OAI21_X2 U11771 ( .B1(n18748), .B2(n11437), .A(n11438), .ZN(n21152) );
  OAI21_X2 U11772 ( .B1(n22388), .B2(n26288), .A(n16341), .ZN(n24811) );
  NOR4_X2 U11773 ( .A1(n26303), .A2(n24891), .A3(n24868), .A4(n22422), .ZN(
        n11639) );
  AOI21_X2 U11774 ( .B1(n16359), .B2(n19349), .A(reset), .ZN(n11634) );
  NOR2_X2 U11775 ( .A1(n22417), .A2(n22416), .ZN(n11200) );
  MUX2_X2 U11776 ( .A(n25769), .B(n25770), .S(n25909), .Z(n25768) );
  OR2_X4 U11777 ( .A1(n12658), .A2(n12659), .ZN(n25770) );
  MUX2_X2 U11778 ( .A(n25772), .B(n25773), .S(n25909), .Z(n25771) );
  OR2_X4 U11779 ( .A1(n12736), .A2(n12737), .ZN(n25773) );
  NAND2_X2 U11780 ( .A1(n22421), .A2(n11874), .ZN(n11806) );
  NAND2_X2 U11781 ( .A1(n25959), .A2(n20458), .ZN(n10081) );
  NAND3_X2 U11782 ( .A1(n22421), .A2(n19348), .A3(n11880), .ZN(n11813) );
  NAND3_X2 U11783 ( .A1(n19348), .A2(n24894), .A3(n11880), .ZN(n11809) );
  AOI21_X2 U11784 ( .B1(n27805), .B2(n25958), .A(n26293), .ZN(n23440) );
  AOI21_X2 U11785 ( .B1(n16374), .B2(n11430), .A(n26293), .ZN(n21149) );
  AOI21_X2 U11786 ( .B1(n22381), .B2(n26267), .A(n26293), .ZN(n24818) );
  AOI21_X2 U11787 ( .B1(n22427), .B2(n26343), .A(n26293), .ZN(n24823) );
  OAI21_X2 U11788 ( .B1(xxx__dut__go), .B2(n16365), .A(n11634), .ZN(n22382) );
  OAI21_X2 U11789 ( .B1(n22401), .B2(n13072), .A(n13073), .ZN(n23445) );
  AOI21_X2 U11790 ( .B1(n11634), .B2(n22402), .A(n11400), .ZN(n13072) );
  OAI21_X2 U11791 ( .B1(n22403), .B2(n13076), .A(n13077), .ZN(n23446) );
  OAI21_X2 U11792 ( .B1(n11794), .B2(dut__bvm__enable), .A(n26350), .ZN(n11793) );
  NOR2_X2 U11793 ( .A1(n25954), .A2(n19539), .ZN(n25774) );
  INV_X4 U11794 ( .A(n2369), .ZN(n26207) );
  INV_X4 U11795 ( .A(n2368), .ZN(n26208) );
  INV_X4 U11796 ( .A(n2367), .ZN(n26209) );
  INV_X4 U11797 ( .A(n2366), .ZN(n26210) );
  INV_X4 U11798 ( .A(n2365), .ZN(n26211) );
  INV_X4 U11799 ( .A(n2364), .ZN(n26212) );
  INV_X4 U11800 ( .A(n2363), .ZN(n26213) );
  INV_X4 U11801 ( .A(n2362), .ZN(n26214) );
  INV_X4 U11802 ( .A(n2361), .ZN(n26215) );
  INV_X4 U11803 ( .A(n2360), .ZN(n26216) );
  INV_X4 U11804 ( .A(n2359), .ZN(n26217) );
  INV_X4 U11805 ( .A(n2358), .ZN(n26218) );
  INV_X4 U11806 ( .A(n2357), .ZN(n26219) );
  INV_X4 U11807 ( .A(n2356), .ZN(n26220) );
  INV_X4 U11808 ( .A(n2355), .ZN(n26221) );
  INV_X4 U11809 ( .A(n2385), .ZN(n26192) );
  INV_X4 U11810 ( .A(n2384), .ZN(n26193) );
  INV_X4 U11811 ( .A(n2383), .ZN(n26194) );
  INV_X4 U11812 ( .A(n2382), .ZN(n26195) );
  INV_X4 U11813 ( .A(n2381), .ZN(n26196) );
  INV_X4 U11814 ( .A(n2380), .ZN(n26197) );
  INV_X4 U11815 ( .A(n2379), .ZN(n26198) );
  INV_X4 U11816 ( .A(n2378), .ZN(n26199) );
  INV_X4 U11817 ( .A(n2377), .ZN(n26200) );
  INV_X4 U11818 ( .A(n2376), .ZN(n26201) );
  INV_X4 U11819 ( .A(n2375), .ZN(n26202) );
  INV_X4 U11820 ( .A(n2374), .ZN(n26203) );
  INV_X4 U11821 ( .A(n2373), .ZN(n26204) );
  INV_X4 U11822 ( .A(n2372), .ZN(n26205) );
  INV_X4 U11823 ( .A(n2371), .ZN(n26206) );
  INV_X4 U11824 ( .A(n2401), .ZN(n26252) );
  INV_X4 U11825 ( .A(n2400), .ZN(n26253) );
  INV_X4 U11826 ( .A(n2399), .ZN(n26254) );
  INV_X4 U11827 ( .A(n2398), .ZN(n26255) );
  INV_X4 U11828 ( .A(n2397), .ZN(n26256) );
  INV_X4 U11829 ( .A(n2396), .ZN(n26257) );
  INV_X4 U11830 ( .A(n2395), .ZN(n26258) );
  INV_X4 U11831 ( .A(n2394), .ZN(n26259) );
  INV_X4 U11832 ( .A(n2393), .ZN(n26260) );
  INV_X4 U11833 ( .A(n2392), .ZN(n26261) );
  INV_X4 U11834 ( .A(n2391), .ZN(n26262) );
  INV_X4 U11835 ( .A(n2390), .ZN(n26263) );
  INV_X4 U11836 ( .A(n2389), .ZN(n26264) );
  INV_X4 U11837 ( .A(n2388), .ZN(n26265) );
  INV_X4 U11838 ( .A(n2387), .ZN(n26266) );
  INV_X4 U11839 ( .A(n2353), .ZN(n26237) );
  INV_X4 U11840 ( .A(n2352), .ZN(n26238) );
  INV_X4 U11841 ( .A(n2351), .ZN(n26239) );
  INV_X4 U11842 ( .A(n2350), .ZN(n26240) );
  INV_X4 U11843 ( .A(n2349), .ZN(n26241) );
  INV_X4 U11844 ( .A(n2348), .ZN(n26242) );
  INV_X4 U11845 ( .A(n2347), .ZN(n26243) );
  INV_X4 U11846 ( .A(n2346), .ZN(n26244) );
  INV_X4 U11847 ( .A(n2345), .ZN(n26245) );
  INV_X4 U11848 ( .A(n2344), .ZN(n26246) );
  INV_X4 U11849 ( .A(n2343), .ZN(n26247) );
  INV_X4 U11850 ( .A(n2342), .ZN(n26248) );
  INV_X4 U11851 ( .A(n2341), .ZN(n26249) );
  INV_X4 U11852 ( .A(n2340), .ZN(n26250) );
  INV_X4 U11853 ( .A(n2339), .ZN(n26251) );
  XNOR2_X2 U11854 ( .A(add_1445_B_7_), .B(n25775), .ZN(U4_DATA1_7) );
  NAND2_X2 U11855 ( .A1(add_1445_B_7_), .A2(add_1445_B_6_), .ZN(n25776) );
  INV_X4 U11856 ( .A(n25776), .ZN(add_1445_carry_8_) );
  XNOR2_X2 U11857 ( .A(add_1445_B_8_), .B(n25776), .ZN(U4_DATA1_8) );
  NAND2_X2 U11858 ( .A1(add_1445_B_8_), .A2(add_1445_carry_8_), .ZN(n25777) );
  XNOR2_X2 U11859 ( .A(add_1445_B_9_), .B(n25777), .ZN(U4_DATA1_9) );
  AND3_X4 U11860 ( .A1(n16216), .A2(n24832), .A3(n22386), .ZN(n25781) );
  AND3_X4 U11861 ( .A1(n22392), .A2(add_180_A_0_), .A3(n25250), .ZN(n12786) );
  AND3_X4 U11862 ( .A1(n22394), .A2(add_180_A_2_), .A3(n25250), .ZN(n12788) );
  AND2_X4 U11863 ( .A1(n16115), .A2(n13032), .ZN(n11501) );
  AND2_X4 U11864 ( .A1(n16115), .A2(n26516), .ZN(n11510) );
  AND2_X4 U11865 ( .A1(n16115), .A2(n26512), .ZN(n11519) );
  AND2_X4 U11866 ( .A1(n16115), .A2(n12889), .ZN(n11528) );
  AND2_X4 U11867 ( .A1(n15977), .A2(n13032), .ZN(n11537) );
  AND2_X4 U11868 ( .A1(n15977), .A2(n26516), .ZN(n11546) );
  AND2_X4 U11869 ( .A1(n15977), .A2(n26512), .ZN(n11555) );
  AND2_X4 U11870 ( .A1(n15977), .A2(n12889), .ZN(n11564) );
  AND2_X4 U11871 ( .A1(n15823), .A2(n13032), .ZN(n11573) );
  AND2_X4 U11872 ( .A1(n15823), .A2(n26516), .ZN(n11582) );
  AND2_X4 U11873 ( .A1(n15823), .A2(n26512), .ZN(n11591) );
  AND2_X4 U11874 ( .A1(n15823), .A2(n12889), .ZN(n11600) );
  AND2_X4 U11875 ( .A1(n13032), .A2(n15606), .ZN(n11419) );
  AND2_X4 U11876 ( .A1(n26516), .A2(n15606), .ZN(n11609) );
  AND2_X4 U11877 ( .A1(n26512), .A2(n15606), .ZN(n11618) );
  AND2_X4 U11878 ( .A1(n12889), .A2(n15606), .ZN(n11627) );
  AND2_X4 U11879 ( .A1(n15526), .A2(n22392), .ZN(n12803) );
  AND2_X4 U11880 ( .A1(n15526), .A2(add_180_A_2_), .ZN(n12811) );
  AND2_X4 U11881 ( .A1(n11794), .A2(n13032), .ZN(n11480) );
  AND2_X2 U11882 ( .A1(n26516), .A2(n11794), .ZN(n11471) );
  AND2_X2 U11883 ( .A1(n26512), .A2(n11794), .ZN(n11462) );
  AND2_X2 U11884 ( .A1(n12889), .A2(n11794), .ZN(n11453) );
  AND2_X4 U11885 ( .A1(n12811), .A2(n12790), .ZN(n12219) );
  AND2_X4 U11886 ( .A1(n12812), .A2(n12790), .ZN(n12221) );
  AND2_X4 U11887 ( .A1(n27799), .A2(n12789), .ZN(n12212) );
  AND2_X4 U11888 ( .A1(n12813), .A2(n12789), .ZN(n12213) );
  AND2_X4 U11889 ( .A1(n12811), .A2(n12791), .ZN(n12203) );
  AND2_X4 U11890 ( .A1(n12812), .A2(n12791), .ZN(n12205) );
  AND2_X4 U11891 ( .A1(n12813), .A2(n12787), .ZN(n12196) );
  AND2_X4 U11892 ( .A1(n12788), .A2(n12787), .ZN(n12197) );
  AND2_X4 U11893 ( .A1(n12803), .A2(n12789), .ZN(n12185) );
  AND2_X4 U11894 ( .A1(n12803), .A2(n12790), .ZN(n12186) );
  AND2_X4 U11895 ( .A1(n12799), .A2(n12789), .ZN(n12177) );
  AND2_X4 U11896 ( .A1(n12799), .A2(n12790), .ZN(n12178) );
  AND2_X4 U11897 ( .A1(n27800), .A2(n12791), .ZN(n12170) );
  AND2_X4 U11898 ( .A1(n27800), .A2(n12789), .ZN(n12172) );
  AND2_X4 U11899 ( .A1(n12786), .A2(n12791), .ZN(n12160) );
  AND2_X4 U11900 ( .A1(n12786), .A2(n12789), .ZN(n12162) );
  AND2_X4 U11901 ( .A1(n11275), .A2(n25247), .ZN(n10207) );
  AND2_X4 U11902 ( .A1(n11276), .A2(n25247), .ZN(n10208) );
  AND2_X4 U11903 ( .A1(n11275), .A2(n11196), .ZN(n10200) );
  AND2_X4 U11904 ( .A1(n11276), .A2(n11196), .ZN(n10201) );
  AND2_X4 U11905 ( .A1(n25247), .A2(n11265), .ZN(n10193) );
  AND2_X4 U11906 ( .A1(n25247), .A2(n11266), .ZN(n10194) );
  AND2_X4 U11907 ( .A1(n11200), .A2(n11265), .ZN(n10186) );
  AND2_X4 U11908 ( .A1(n11266), .A2(n11200), .ZN(n10187) );
  AND2_X4 U11909 ( .A1(n11227), .A2(n25247), .ZN(n10174) );
  AND2_X4 U11910 ( .A1(n11221), .A2(n25247), .ZN(n10175) );
  AND2_X4 U11911 ( .A1(n11227), .A2(n11196), .ZN(n10167) );
  AND2_X4 U11912 ( .A1(n11225), .A2(n11195), .ZN(n10168) );
  AND2_X4 U11913 ( .A1(n11244), .A2(n25247), .ZN(n10160) );
  AND2_X4 U11914 ( .A1(n11245), .A2(n25247), .ZN(n10161) );
  AND2_X4 U11915 ( .A1(n11244), .A2(n11196), .ZN(n10153) );
  AND2_X4 U11916 ( .A1(n11245), .A2(n11196), .ZN(n10154) );
  AND2_X4 U11917 ( .A1(n11231), .A2(n11196), .ZN(n10142) );
  AND2_X4 U11918 ( .A1(n11226), .A2(n11200), .ZN(n10144) );
  AND2_X4 U11919 ( .A1(n11231), .A2(n11195), .ZN(n10135) );
  AND2_X4 U11920 ( .A1(n11226), .A2(n11196), .ZN(n10137) );
  AND2_X4 U11921 ( .A1(n11220), .A2(n11196), .ZN(n10128) );
  AND2_X4 U11922 ( .A1(n11227), .A2(n11200), .ZN(n10130) );
  AND2_X4 U11923 ( .A1(n11220), .A2(n11195), .ZN(n10121) );
  AND2_X4 U11924 ( .A1(n11221), .A2(n11196), .ZN(n10123) );
  AND2_X4 U11925 ( .A1(n11207), .A2(n11200), .ZN(n10111) );
  AND2_X4 U11926 ( .A1(n11207), .A2(n11195), .ZN(n10104) );
  AND2_X4 U11927 ( .A1(n24886), .A2(n11196), .ZN(n10106) );
  AND2_X4 U11928 ( .A1(n11192), .A2(n11196), .ZN(n10097) );
  AND2_X4 U11929 ( .A1(n11194), .A2(n11200), .ZN(n10099) );
  AND2_X4 U11930 ( .A1(n11192), .A2(n11195), .ZN(n10090) );
  AND2_X4 U11931 ( .A1(n11194), .A2(n11196), .ZN(n10092) );
  NAND2_X2 U11932 ( .A1(n26135), .A2(n26137), .ZN(n11283) );
  MUX2_X2 U11933 ( .A(n20524), .B(n26134), .S(n25959), .Z(n25985) );
  INV_X4 U11934 ( .A(n25985), .ZN(n20556) );
  INV_X4 U11935 ( .A(n25986), .ZN(n20557) );
  MUX2_X2 U11936 ( .A(n20526), .B(n26132), .S(n25959), .Z(n25987) );
  INV_X4 U11937 ( .A(n25987), .ZN(n20558) );
  MUX2_X2 U11938 ( .A(n25778), .B(n26131), .S(n25959), .Z(n25988) );
  INV_X4 U11939 ( .A(n25988), .ZN(n20559) );
  NOR4_X2 U11940 ( .A1(n11181), .A2(n11182), .A3(n11183), .A4(n11184), .ZN(
        n25989) );
  MUX2_X2 U11941 ( .A(n20523), .B(n25989), .S(n26130), .Z(n25990) );
  INV_X4 U11942 ( .A(n25990), .ZN(n20555) );
  NOR4_X2 U11943 ( .A1(n11112), .A2(n11113), .A3(n11114), .A4(n11115), .ZN(
        n25991) );
  INV_X4 U11944 ( .A(n25992), .ZN(n20554) );
  NOR4_X2 U11945 ( .A1(n11043), .A2(n11044), .A3(n11045), .A4(n11046), .ZN(
        n25993) );
  MUX2_X2 U11946 ( .A(n20392), .B(n25993), .S(n26130), .Z(n25994) );
  INV_X4 U11947 ( .A(n25994), .ZN(n20553) );
  NOR4_X2 U11948 ( .A1(n10974), .A2(n10975), .A3(n10976), .A4(n10977), .ZN(
        n25995) );
  MUX2_X2 U11949 ( .A(n25750), .B(n25995), .S(n26130), .Z(n25996) );
  INV_X4 U11950 ( .A(n25996), .ZN(n20552) );
  NOR4_X2 U11951 ( .A1(n10905), .A2(n10906), .A3(n10907), .A4(n10908), .ZN(
        n25997) );
  MUX2_X2 U11952 ( .A(n20262), .B(n25997), .S(n26130), .Z(n25998) );
  INV_X4 U11953 ( .A(n25998), .ZN(n20551) );
  NOR4_X2 U11954 ( .A1(n10836), .A2(n10837), .A3(n10838), .A4(n10839), .ZN(
        n25999) );
  INV_X4 U11955 ( .A(n26000), .ZN(n20550) );
  NOR2_X2 U11957 ( .A1(n12775), .A2(n12776), .ZN(n26001) );
  MUX2_X2 U11958 ( .A(n18792), .B(n26001), .S(n25909), .Z(n26002) );
  INV_X4 U11959 ( .A(n26002), .ZN(n23103) );
  NOR2_X2 U11960 ( .A1(n12697), .A2(n12698), .ZN(n26003) );
  MUX2_X2 U11961 ( .A(n18866), .B(n26003), .S(n25909), .Z(n26004) );
  INV_X4 U11962 ( .A(n26004), .ZN(n23101) );
  NOR2_X2 U11963 ( .A1(n12619), .A2(n12620), .ZN(n26005) );
  MUX2_X2 U11964 ( .A(n18940), .B(n26005), .S(n25909), .Z(n26006) );
  INV_X4 U11965 ( .A(n26006), .ZN(n23099) );
  NOR2_X2 U11966 ( .A1(n12580), .A2(n12581), .ZN(n26007) );
  MUX2_X2 U11967 ( .A(n18977), .B(n26007), .S(n25909), .Z(n26008) );
  INV_X4 U11968 ( .A(n26008), .ZN(n23098) );
  NOR2_X2 U11969 ( .A1(n12541), .A2(n12542), .ZN(n26009) );
  MUX2_X2 U11970 ( .A(n19014), .B(n26009), .S(n25909), .Z(n26010) );
  INV_X4 U11971 ( .A(n26010), .ZN(n23097) );
  NOR2_X2 U11972 ( .A1(n12502), .A2(n12503), .ZN(n26011) );
  MUX2_X2 U11973 ( .A(n25976), .B(n26011), .S(n25909), .Z(n26012) );
  NOR2_X2 U11974 ( .A1(n12463), .A2(n12464), .ZN(n26013) );
  MUX2_X2 U11975 ( .A(n19088), .B(n26013), .S(n25909), .Z(n26014) );
  INV_X4 U11976 ( .A(n26014), .ZN(n23095) );
  NOR2_X2 U11977 ( .A1(n12424), .A2(n12425), .ZN(n26015) );
  MUX2_X2 U11978 ( .A(n25973), .B(n26015), .S(n25909), .Z(n26016) );
  INV_X4 U11979 ( .A(n26016), .ZN(n23094) );
  NOR2_X2 U11980 ( .A1(n12385), .A2(n12386), .ZN(n26017) );
  MUX2_X2 U11981 ( .A(n25971), .B(n26017), .S(n25907), .Z(n26018) );
  INV_X4 U11982 ( .A(n26018), .ZN(n23093) );
  NOR2_X2 U11983 ( .A1(n12346), .A2(n12347), .ZN(n26019) );
  MUX2_X2 U11984 ( .A(n25969), .B(n26019), .S(n25909), .Z(n26020) );
  INV_X4 U11985 ( .A(n26020), .ZN(n23092) );
  NOR2_X2 U11986 ( .A1(n14911), .A2(n14912), .ZN(n26021) );
  MUX2_X2 U11987 ( .A(n16966), .B(n26021), .S(n25909), .Z(n26022) );
  INV_X4 U11988 ( .A(n26022), .ZN(n23500) );
  NOR2_X2 U11989 ( .A1(n14948), .A2(n14949), .ZN(n26023) );
  INV_X4 U11990 ( .A(n26024), .ZN(n23501) );
  NOR2_X2 U11991 ( .A1(n14985), .A2(n14986), .ZN(n26025) );
  MUX2_X2 U11992 ( .A(n16892), .B(n26025), .S(n25907), .Z(n26026) );
  INV_X4 U11993 ( .A(n26026), .ZN(n23502) );
  NOR2_X2 U11994 ( .A1(n15022), .A2(n15023), .ZN(n26027) );
  MUX2_X2 U11995 ( .A(n25740), .B(n26027), .S(n25907), .Z(n26028) );
  INV_X4 U11996 ( .A(n26028), .ZN(n23503) );
  NOR2_X2 U11997 ( .A1(n15059), .A2(n15060), .ZN(n26029) );
  MUX2_X2 U11998 ( .A(n16818), .B(n26029), .S(n25907), .Z(n26030) );
  INV_X4 U11999 ( .A(n26030), .ZN(n23504) );
  NOR2_X2 U12000 ( .A1(n15096), .A2(n15097), .ZN(n26031) );
  INV_X4 U12001 ( .A(n26032), .ZN(n23505) );
  NOR2_X2 U12002 ( .A1(n14319), .A2(n14320), .ZN(n26033) );
  MUX2_X2 U12003 ( .A(n17558), .B(n26033), .S(n25909), .Z(n26034) );
  INV_X4 U12004 ( .A(n26034), .ZN(n23484) );
  NOR2_X2 U12005 ( .A1(n14356), .A2(n14357), .ZN(n26035) );
  MUX2_X2 U12006 ( .A(n17521), .B(n26035), .S(n25909), .Z(n26036) );
  INV_X4 U12007 ( .A(n26036), .ZN(n23485) );
  NOR2_X2 U12008 ( .A1(n14393), .A2(n14394), .ZN(n26037) );
  MUX2_X2 U12009 ( .A(n17484), .B(n26037), .S(n25907), .Z(n26038) );
  INV_X4 U12010 ( .A(n26038), .ZN(n23486) );
  NOR2_X2 U12011 ( .A1(n14430), .A2(n14431), .ZN(n26039) );
  MUX2_X2 U12012 ( .A(n17447), .B(n26039), .S(n25909), .Z(n26040) );
  INV_X4 U12013 ( .A(n26040), .ZN(n23487) );
  NOR2_X2 U12014 ( .A1(n14467), .A2(n14468), .ZN(n26041) );
  MUX2_X2 U12015 ( .A(n17410), .B(n26041), .S(n25909), .Z(n26042) );
  INV_X4 U12016 ( .A(n26042), .ZN(n23488) );
  NOR2_X2 U12017 ( .A1(n14504), .A2(n14505), .ZN(n26043) );
  MUX2_X2 U12018 ( .A(n17373), .B(n26043), .S(n25907), .Z(n26044) );
  INV_X4 U12019 ( .A(n26044), .ZN(n23489) );
  NOR2_X2 U12020 ( .A1(n14541), .A2(n14542), .ZN(n26045) );
  MUX2_X2 U12021 ( .A(n17336), .B(n26045), .S(n25907), .Z(n26046) );
  INV_X4 U12022 ( .A(n26046), .ZN(n23490) );
  NOR2_X2 U12023 ( .A1(n14578), .A2(n14579), .ZN(n26047) );
  MUX2_X2 U12024 ( .A(n17299), .B(n26047), .S(n25907), .Z(n26048) );
  INV_X4 U12025 ( .A(n26048), .ZN(n23491) );
  NOR2_X2 U12026 ( .A1(n14615), .A2(n14616), .ZN(n26049) );
  MUX2_X2 U12027 ( .A(n17262), .B(n26049), .S(n25907), .Z(n26050) );
  INV_X4 U12028 ( .A(n26050), .ZN(n23492) );
  NOR2_X2 U12029 ( .A1(n14652), .A2(n14653), .ZN(n26051) );
  MUX2_X2 U12030 ( .A(n17225), .B(n26051), .S(n25907), .Z(n26052) );
  INV_X4 U12031 ( .A(n26052), .ZN(n23493) );
  NOR2_X2 U12032 ( .A1(n14689), .A2(n14690), .ZN(n26053) );
  MUX2_X2 U12033 ( .A(n17188), .B(n26053), .S(n25907), .Z(n26054) );
  INV_X4 U12034 ( .A(n26054), .ZN(n23494) );
  NOR2_X2 U12035 ( .A1(n14726), .A2(n14727), .ZN(n26055) );
  MUX2_X2 U12036 ( .A(n17151), .B(n26055), .S(n25907), .Z(n26056) );
  INV_X4 U12037 ( .A(n26056), .ZN(n23495) );
  NOR2_X2 U12038 ( .A1(n13727), .A2(n13728), .ZN(n26057) );
  MUX2_X2 U12039 ( .A(n18150), .B(n26057), .S(n25907), .Z(n26058) );
  INV_X4 U12040 ( .A(n26058), .ZN(n23468) );
  NOR2_X2 U12041 ( .A1(n13764), .A2(n13765), .ZN(n26059) );
  MUX2_X2 U12042 ( .A(n18113), .B(n26059), .S(n25907), .Z(n26060) );
  INV_X4 U12043 ( .A(n26060), .ZN(n23469) );
  NOR2_X2 U12044 ( .A1(n13801), .A2(n13802), .ZN(n26061) );
  MUX2_X2 U12045 ( .A(n18076), .B(n26061), .S(n25907), .Z(n26062) );
  INV_X4 U12046 ( .A(n26062), .ZN(n23470) );
  NOR2_X2 U12047 ( .A1(n13838), .A2(n13839), .ZN(n26063) );
  MUX2_X2 U12048 ( .A(n18039), .B(n26063), .S(n25907), .Z(n26064) );
  INV_X4 U12049 ( .A(n26064), .ZN(n23471) );
  NOR2_X2 U12050 ( .A1(n13875), .A2(n13876), .ZN(n26065) );
  MUX2_X2 U12051 ( .A(n18002), .B(n26065), .S(n25907), .Z(n26066) );
  INV_X4 U12052 ( .A(n26066), .ZN(n23472) );
  NOR2_X2 U12053 ( .A1(n13912), .A2(n13913), .ZN(n26067) );
  MUX2_X2 U12054 ( .A(n17965), .B(n26067), .S(n25907), .Z(n26068) );
  INV_X4 U12055 ( .A(n26068), .ZN(n23473) );
  NOR2_X2 U12056 ( .A1(n13949), .A2(n13950), .ZN(n26069) );
  MUX2_X2 U12057 ( .A(n17928), .B(n26069), .S(n25907), .Z(n26070) );
  INV_X4 U12058 ( .A(n26070), .ZN(n23474) );
  NOR2_X2 U12059 ( .A1(n13986), .A2(n13987), .ZN(n26071) );
  MUX2_X2 U12060 ( .A(n17891), .B(n26071), .S(n25907), .Z(n26072) );
  INV_X4 U12061 ( .A(n26072), .ZN(n23475) );
  NOR2_X2 U12062 ( .A1(n14023), .A2(n14024), .ZN(n26073) );
  MUX2_X2 U12063 ( .A(n17854), .B(n26073), .S(n25907), .Z(n26074) );
  INV_X4 U12064 ( .A(n26074), .ZN(n23476) );
  NOR2_X2 U12065 ( .A1(n14060), .A2(n14061), .ZN(n26075) );
  MUX2_X2 U12066 ( .A(n17817), .B(n26075), .S(n25909), .Z(n26076) );
  INV_X4 U12067 ( .A(n26076), .ZN(n23477) );
  NOR2_X2 U12068 ( .A1(n14097), .A2(n14098), .ZN(n26077) );
  MUX2_X2 U12069 ( .A(n17780), .B(n26077), .S(n25909), .Z(n26078) );
  INV_X4 U12070 ( .A(n26078), .ZN(n23478) );
  NOR2_X2 U12071 ( .A1(n14134), .A2(n14135), .ZN(n26079) );
  MUX2_X2 U12072 ( .A(n17743), .B(n26079), .S(n25909), .Z(n26080) );
  INV_X4 U12073 ( .A(n26080), .ZN(n23479) );
  NOR2_X2 U12074 ( .A1(n13099), .A2(n13100), .ZN(n26081) );
  MUX2_X2 U12075 ( .A(n18742), .B(n26081), .S(n25909), .Z(n26082) );
  INV_X4 U12076 ( .A(n26082), .ZN(n23452) );
  NOR2_X2 U12077 ( .A1(n13172), .A2(n13173), .ZN(n26083) );
  MUX2_X2 U12078 ( .A(n18705), .B(n26083), .S(n25909), .Z(n26084) );
  INV_X4 U12079 ( .A(n26084), .ZN(n23453) );
  NOR2_X2 U12080 ( .A1(n13209), .A2(n13210), .ZN(n26085) );
  MUX2_X2 U12081 ( .A(n18668), .B(n26085), .S(n25909), .Z(n26086) );
  INV_X4 U12082 ( .A(n26086), .ZN(n23454) );
  NOR2_X2 U12083 ( .A1(n13246), .A2(n13247), .ZN(n26087) );
  MUX2_X2 U12084 ( .A(n18631), .B(n26087), .S(n25909), .Z(n26088) );
  INV_X4 U12085 ( .A(n26088), .ZN(n23455) );
  NOR2_X2 U12086 ( .A1(n13283), .A2(n13284), .ZN(n26089) );
  MUX2_X2 U12087 ( .A(n18594), .B(n26089), .S(n25909), .Z(n26090) );
  INV_X4 U12088 ( .A(n26090), .ZN(n23456) );
  NOR2_X2 U12089 ( .A1(n13320), .A2(n13321), .ZN(n26091) );
  MUX2_X2 U12090 ( .A(n18557), .B(n26091), .S(n25909), .Z(n26092) );
  INV_X4 U12091 ( .A(n26092), .ZN(n23457) );
  NOR2_X2 U12092 ( .A1(n13357), .A2(n13358), .ZN(n26093) );
  MUX2_X2 U12093 ( .A(n18520), .B(n26093), .S(n25909), .Z(n26094) );
  INV_X4 U12094 ( .A(n26094), .ZN(n23458) );
  NOR2_X2 U12095 ( .A1(n13394), .A2(n13395), .ZN(n26095) );
  MUX2_X2 U12096 ( .A(n18483), .B(n26095), .S(n25909), .Z(n26096) );
  INV_X4 U12097 ( .A(n26096), .ZN(n23459) );
  NOR2_X2 U12098 ( .A1(n13431), .A2(n13432), .ZN(n26097) );
  MUX2_X2 U12099 ( .A(n18446), .B(n26097), .S(n25909), .Z(n26098) );
  INV_X4 U12100 ( .A(n26098), .ZN(n23460) );
  NOR2_X2 U12101 ( .A1(n13468), .A2(n13469), .ZN(n26099) );
  MUX2_X2 U12102 ( .A(n18409), .B(n26099), .S(n25909), .Z(n26100) );
  INV_X4 U12103 ( .A(n26100), .ZN(n23461) );
  NOR2_X2 U12104 ( .A1(n13505), .A2(n13506), .ZN(n26101) );
  MUX2_X2 U12105 ( .A(n18372), .B(n26101), .S(n25909), .Z(n26102) );
  INV_X4 U12106 ( .A(n26102), .ZN(n23462) );
  NOR2_X2 U12107 ( .A1(n13542), .A2(n13543), .ZN(n26103) );
  MUX2_X2 U12108 ( .A(n18335), .B(n26103), .S(n25909), .Z(n26104) );
  INV_X4 U12109 ( .A(n26104), .ZN(n23463) );
  NAND3_X2 U12110 ( .A1(n19348), .A2(n24894), .A3(n25255), .ZN(n26105) );
  NAND2_X2 U12111 ( .A1(n26105), .A2(n26139), .ZN(n26107) );
  INV_X4 U12112 ( .A(n26107), .ZN(n26106) );
  NAND2_X2 U12113 ( .A1(n26106), .A2(n11634), .ZN(n26110) );
  NOR2_X2 U12114 ( .A1(n26296), .A2(n26110), .ZN(n26109) );
  NAND3_X2 U12115 ( .A1(n13043), .A2(n11634), .A3(n26107), .ZN(n26108) );
  NAND2_X2 U12116 ( .A1(n26108), .A2(n11441), .ZN(n26115) );
  MUX2_X2 U12117 ( .A(n26109), .B(n26115), .S(n19348), .Z(n23433) );
  INV_X4 U12118 ( .A(n26115), .ZN(n26112) );
  INV_X4 U12119 ( .A(n26110), .ZN(n26116) );
  NAND2_X2 U12120 ( .A1(n26116), .A2(n26129), .ZN(n26111) );
  NAND2_X2 U12121 ( .A1(n26112), .A2(n26111), .ZN(n26114) );
  NAND3_X2 U12122 ( .A1(n26116), .A2(n19348), .A3(n11441), .ZN(n26117) );
  INV_X4 U12123 ( .A(n26117), .ZN(n26113) );
  MUX2_X2 U12124 ( .A(n26114), .B(n26113), .S(n22421), .Z(n23432) );
  NOR2_X2 U12125 ( .A1(n26116), .A2(n26115), .ZN(n26118) );
  OAI22_X2 U12126 ( .A1(n22420), .A2(n26118), .B1(n22421), .B2(n26117), .ZN(
        n23431) );
  INV_X4 U12127 ( .A(n16364), .ZN(n26120) );
  INV_X4 U12128 ( .A(n16358), .ZN(n26119) );
  MUX2_X2 U12129 ( .A(n26120), .B(n26119), .S(n22424), .Z(n24822) );
  NOR2_X2 U12130 ( .A1(n22424), .A2(n16358), .ZN(n26121) );
  MUX2_X2 U12131 ( .A(n16361), .B(n26121), .S(n22423), .Z(n24821) );
  NAND3_X2 U12132 ( .A1(n22422), .A2(n24891), .A3(n24868), .ZN(n11788) );
  NAND2_X2 U12133 ( .A1(n22385), .A2(n24833), .ZN(n16354) );
  INV_X4 U12134 ( .A(n16348), .ZN(n26122) );
  NAND4_X2 U12135 ( .A1(n22384), .A2(n24833), .A3(n25400), .A4(n26122), .ZN(
        n16351) );
  NAND2_X2 U12136 ( .A1(n22390), .A2(n25256), .ZN(n26514) );
  NAND2_X2 U12137 ( .A1(n22389), .A2(n25254), .ZN(n16192) );
  INV_X4 U12138 ( .A(n26514), .ZN(n12889) );
  INV_X4 U12139 ( .A(n16192), .ZN(n26512) );
  NAND2_X2 U12140 ( .A1(n22393), .A2(add_180_A_0_), .ZN(n15546) );
  INV_X4 U12141 ( .A(n15538), .ZN(n26285) );
  INV_X4 U12142 ( .A(n15539), .ZN(n26123) );
  NAND4_X2 U12143 ( .A1(add_180_A_0_), .A2(add_180_A_1_), .A3(n22392), .A4(
        n26123), .ZN(n15543) );
  NAND2_X2 U12144 ( .A1(n15513), .A2(n22396), .ZN(n15534) );
  NAND2_X2 U12145 ( .A1(n13075), .A2(n22406), .ZN(n13092) );
  NAND2_X2 U12146 ( .A1(n22404), .A2(n25104), .ZN(n13088) );
  INV_X4 U12147 ( .A(n13084), .ZN(n26124) );
  NAND4_X2 U12148 ( .A1(n25104), .A2(n26136), .A3(n25401), .A4(n26124), .ZN(
        n13083) );
  INV_X4 U12149 ( .A(n13078), .ZN(n26138) );
  NAND4_X2 U12150 ( .A1(n22403), .A2(n13075), .A3(n11634), .A4(n26138), .ZN(
        n13077) );
  INV_X4 U12151 ( .A(n11399), .ZN(n26125) );
  NAND3_X2 U12152 ( .A1(n24887), .A2(n22401), .A3(n26125), .ZN(n13073) );
  NAND2_X2 U12153 ( .A1(n24896), .A2(n24887), .ZN(n13071) );
  INV_X4 U12154 ( .A(add_283_carry[5]), .ZN(n26126) );
  NAND3_X2 U12155 ( .A1(n11878), .A2(n11634), .A3(n26126), .ZN(n26127) );
  NAND2_X2 U12156 ( .A1(n26127), .A2(n13054), .ZN(n26128) );
  NAND2_X2 U12157 ( .A1(add_283_A_5_), .A2(n26128), .ZN(n13045) );
  INV_X4 U12158 ( .A(n11400), .ZN(n26281) );
  INV_X4 U12159 ( .A(n[618]), .ZN(n26222) );
  INV_X4 U12160 ( .A(n[617]), .ZN(n26223) );
  INV_X4 U12161 ( .A(n[616]), .ZN(n26224) );
  INV_X4 U12162 ( .A(n[615]), .ZN(n26225) );
  INV_X4 U12163 ( .A(n[614]), .ZN(n26226) );
  INV_X4 U12164 ( .A(n[613]), .ZN(n26227) );
  INV_X4 U12165 ( .A(n[612]), .ZN(n26228) );
  INV_X4 U12166 ( .A(n[611]), .ZN(n26229) );
  INV_X4 U12167 ( .A(n[610]), .ZN(n26230) );
  INV_X4 U12168 ( .A(n[609]), .ZN(n26231) );
  INV_X4 U12169 ( .A(n[608]), .ZN(n26232) );
  INV_X4 U12170 ( .A(n[607]), .ZN(n26233) );
  INV_X4 U12171 ( .A(n[606]), .ZN(n26234) );
  INV_X4 U12172 ( .A(n[605]), .ZN(n26235) );
  INV_X4 U12173 ( .A(n[604]), .ZN(n26236) );
  INV_X4 U12174 ( .A(xxx__dut__go), .ZN(n26267) );
  INV_X4 U12175 ( .A(n13059), .ZN(n26280) );
  INV_X4 U12176 ( .A(n13086), .ZN(n26282) );
  INV_X4 U12177 ( .A(n13085), .ZN(n26283) );
  INV_X4 U12178 ( .A(n15541), .ZN(n26284) );
  INV_X4 U12179 ( .A(n15535), .ZN(n26286) );
  INV_X4 U12180 ( .A(n15537), .ZN(n26287) );
  INV_X4 U12181 ( .A(n16343), .ZN(n26288) );
  INV_X4 U12182 ( .A(n16352), .ZN(n26289) );
  INV_X4 U12183 ( .A(n16347), .ZN(n26290) );
  INV_X4 U12184 ( .A(n16342), .ZN(n26291) );
  INV_X4 U12185 ( .A(n16346), .ZN(n26292) );
  INV_X4 U12186 ( .A(n13095), .ZN(n26294) );
  INV_X4 U12187 ( .A(n13075), .ZN(n26295) );
  INV_X4 U12188 ( .A(n11441), .ZN(n26296) );
  INV_X4 U12189 ( .A(n13050), .ZN(n26297) );
  INV_X4 U12190 ( .A(n13051), .ZN(n26298) );
  INV_X4 U12191 ( .A(n13052), .ZN(n26299) );
  INV_X4 U12192 ( .A(n13053), .ZN(n26300) );
  INV_X4 U12193 ( .A(n13054), .ZN(n26301) );
  INV_X4 U12194 ( .A(n13055), .ZN(n26302) );
  INV_X4 U12195 ( .A(n11434), .ZN(n26304) );
  INV_X4 U12196 ( .A(n16359), .ZN(n26305) );
  INV_X4 U12197 ( .A(n13093), .ZN(n26350) );
  INV_X4 U12198 ( .A(n16179), .ZN(n26459) );
  INV_X4 U12199 ( .A(n11487), .ZN(n26460) );
  INV_X4 U12200 ( .A(n11496), .ZN(n26461) );
  INV_X4 U12201 ( .A(n16196), .ZN(n26498) );
  INV_X4 U12202 ( .A(n11490), .ZN(n26499) );
  INV_X4 U12203 ( .A(n16178), .ZN(n26501) );
  INV_X4 U12204 ( .A(n16207), .ZN(n26503) );
  INV_X4 U12205 ( .A(n12847), .ZN(n26504) );
  INV_X4 U12206 ( .A(n16174), .ZN(n26505) );
  INV_X4 U12207 ( .A(n12978), .ZN(n26507) );
  INV_X4 U12208 ( .A(n12974), .ZN(n26511) );
  INV_X4 U12209 ( .A(n11497), .ZN(n26513) );
  INV_X4 U12210 ( .A(n12975), .ZN(n26515) );
  INV_X4 U12211 ( .A(n16188), .ZN(n26516) );
  INV_X4 U12212 ( .A(n11491), .ZN(n26517) );
  INV_X4 U12213 ( .A(n16191), .ZN(n26518) );
  INV_X4 U12214 ( .A(n15488), .ZN(n27799) );
  INV_X4 U12215 ( .A(n15484), .ZN(n27800) );
  INV_X4 U12216 ( .A(n12826), .ZN(n27801) );
  INV_X4 U12217 ( .A(n15518), .ZN(n27802) );
  INV_X4 U12218 ( .A(n15517), .ZN(n27803) );
  INV_X4 U12219 ( .A(n15514), .ZN(n27804) );
  INV_X4 U12220 ( .A(U8_DATA2_8), .ZN(n27806) );
  INV_X4 U12221 ( .A(U8_DATA2_7), .ZN(n27807) );
  INV_X4 U12222 ( .A(U8_DATA2_6), .ZN(n27808) );
  INV_X4 U12223 ( .A(U8_DATA2_5), .ZN(n27809) );
  INV_X4 U12224 ( .A(U8_DATA2_4), .ZN(n27810) );
  INV_X4 U12225 ( .A(U8_DATA2_3), .ZN(n27811) );
  INV_X4 U12226 ( .A(U8_DATA2_2), .ZN(n27812) );
  INV_X4 U12227 ( .A(U8_DATA2_1), .ZN(n27813) );
  OAI22_X1 U10532 ( .A1(n25950), .A2(n28244), .B1(n26253), .B2(n24845), .ZN(
        n22598) );
  OAI22_X1 U10533 ( .A1(n25950), .A2(n28220), .B1(n26256), .B2(n24845), .ZN(
        n22622) );
  OAI22_X1 U10534 ( .A1(n25951), .A2(n28485), .B1(n26210), .B2(n24845), .ZN(
        n22861) );
  OAI22_X1 U10535 ( .A1(n25951), .A2(n28478), .B1(n26211), .B2(n24845), .ZN(
        n22867) );
  OAI22_X1 U10536 ( .A1(n24846), .A2(n26221), .B1(n20498), .B2(n25956), .ZN(
        n20572) );
  OAI22_X1 U10537 ( .A1(n24846), .A2(n26192), .B1(n19583), .B2(n25956), .ZN(
        n20602) );
  OAI22_X1 U10538 ( .A1(n24846), .A2(n26258), .B1(n25957), .B2(n28205), .ZN(
        n22639) );
  OAI22_X1 U10539 ( .A1(n24846), .A2(n26260), .B1(n25957), .B2(n28189), .ZN(
        n22655) );
  OAI22_X1 U11367 ( .A1(n24846), .A2(n26262), .B1(n25957), .B2(n28173), .ZN(
        n22671) );
  OAI22_X1 U11956 ( .A1(n20519), .A2(n25954), .B1(n26221), .B2(n24864), .ZN(
        n20604) );
  OAI22_X1 U12228 ( .A1(n20453), .A2(n25954), .B1(n26220), .B2(n24864), .ZN(
        n20605) );
  OAI22_X1 U12229 ( .A1(n20388), .A2(n25954), .B1(n26219), .B2(n24864), .ZN(
        n20606) );
  OAI22_X1 U12230 ( .A1(n20323), .A2(n25953), .B1(n26218), .B2(n24864), .ZN(
        n20607) );
  OAI22_X1 U12231 ( .A1(n25953), .A2(n28377), .B1(n26192), .B2(n24864), .ZN(
        n22719) );
  OAI22_X1 U12232 ( .A1(n25953), .A2(n28353), .B1(n26195), .B2(n24864), .ZN(
        n22743) );
  OAI22_X1 U12233 ( .A1(n20512), .A2(n25936), .B1(n26251), .B2(n24889), .ZN(
        n20796) );
  OAI22_X1 U12234 ( .A1(n20446), .A2(n25936), .B1(n26250), .B2(n24889), .ZN(
        n20797) );
  OAI22_X1 U12235 ( .A1(n20381), .A2(n25935), .B1(n26249), .B2(n24889), .ZN(
        n20798) );
  OAI22_X1 U12236 ( .A1(n20316), .A2(n25935), .B1(n26248), .B2(n24889), .ZN(
        n20799) );
  OAI22_X1 U12237 ( .A1(n25935), .A2(n28248), .B1(n26252), .B2(n24889), .ZN(
        n22586) );
  OAI22_X1 U12238 ( .A1(n25935), .A2(n28240), .B1(n26253), .B2(n24889), .ZN(
        n22594) );
  OAI22_X1 U12239 ( .A1(n20513), .A2(n25915), .B1(n26251), .B2(n24888), .ZN(
        n21020) );
  OAI22_X1 U12240 ( .A1(n20447), .A2(n25915), .B1(n26250), .B2(n24888), .ZN(
        n21021) );
  OAI22_X1 U12241 ( .A1(n20382), .A2(n25914), .B1(n26249), .B2(n24888), .ZN(
        n21022) );
  OAI22_X1 U12242 ( .A1(n20317), .A2(n25914), .B1(n26248), .B2(n24888), .ZN(
        n21023) );
  OAI22_X1 U12243 ( .A1(n25914), .A2(n28247), .B1(n26252), .B2(n24888), .ZN(
        n22585) );
  OAI22_X1 U12244 ( .A1(n25914), .A2(n28239), .B1(n26253), .B2(n24888), .ZN(
        n22593) );
  OAI22_X1 U12245 ( .A1(n20511), .A2(n25948), .B1(n26251), .B2(n24844), .ZN(
        n20668) );
  OAI22_X1 U12246 ( .A1(n20445), .A2(n25948), .B1(n26250), .B2(n24844), .ZN(
        n20669) );
  OAI22_X1 U12247 ( .A1(n20380), .A2(n25947), .B1(n26249), .B2(n24844), .ZN(
        n20670) );
  OAI22_X1 U12248 ( .A1(n20315), .A2(n25947), .B1(n26248), .B2(n24844), .ZN(
        n20671) );
  OAI22_X1 U12249 ( .A1(n25947), .A2(n28249), .B1(n26252), .B2(n24844), .ZN(
        n22587) );
  OAI22_X1 U12250 ( .A1(n25947), .A2(n28241), .B1(n26253), .B2(n24844), .ZN(
        n22595) );
  OAI22_X1 U12251 ( .A1(n20503), .A2(n25945), .B1(n26221), .B2(n24843), .ZN(
        n20700) );
  OAI22_X1 U12252 ( .A1(n20437), .A2(n25945), .B1(n26220), .B2(n24843), .ZN(
        n20701) );
  OAI22_X1 U12253 ( .A1(n20372), .A2(n25944), .B1(n26219), .B2(n24843), .ZN(
        n20702) );
  OAI22_X1 U12254 ( .A1(n20307), .A2(n25944), .B1(n26218), .B2(n24843), .ZN(
        n20703) );
  OAI22_X1 U12255 ( .A1(n25944), .A2(n28373), .B1(n26192), .B2(n24843), .ZN(
        n22715) );
  OAI22_X1 U12256 ( .A1(n25944), .A2(n28365), .B1(n26193), .B2(n24843), .ZN(
        n22723) );
  OAI22_X1 U12257 ( .A1(n20520), .A2(n25942), .B1(n26221), .B2(n24842), .ZN(
        n20732) );
  OAI22_X1 U12258 ( .A1(n20454), .A2(n25942), .B1(n26220), .B2(n24842), .ZN(
        n20733) );
  OAI22_X1 U12259 ( .A1(n20389), .A2(n25941), .B1(n26219), .B2(n24842), .ZN(
        n20734) );
  OAI22_X1 U12260 ( .A1(n20324), .A2(n25941), .B1(n26218), .B2(n24842), .ZN(
        n20735) );
  OAI22_X1 U12261 ( .A1(n25941), .A2(n28375), .B1(n26192), .B2(n24842), .ZN(
        n22717) );
  OAI22_X1 U12262 ( .A1(n25941), .A2(n28367), .B1(n26193), .B2(n24842), .ZN(
        n22725) );
  OAI22_X1 U12263 ( .A1(n20365), .A2(n25938), .B1(n26249), .B2(n24841), .ZN(
        n20766) );
  OAI22_X1 U12264 ( .A1(n20300), .A2(n25938), .B1(n26248), .B2(n24841), .ZN(
        n20767) );
  OAI22_X1 U12265 ( .A1(n20235), .A2(n25938), .B1(n26247), .B2(n24841), .ZN(
        n20768) );
  OAI22_X1 U12266 ( .A1(n20170), .A2(n25938), .B1(n26246), .B2(n24841), .ZN(
        n20769) );
  OAI22_X1 U12267 ( .A1(n20105), .A2(n25938), .B1(n26245), .B2(n24841), .ZN(
        n20770) );
  OAI22_X1 U12268 ( .A1(n20040), .A2(n25938), .B1(n26244), .B2(n24841), .ZN(
        n20771) );
  OAI22_X1 U12269 ( .A1(n20504), .A2(n25933), .B1(n26221), .B2(n24840), .ZN(
        n20828) );
  OAI22_X1 U12270 ( .A1(n20438), .A2(n25933), .B1(n26220), .B2(n24840), .ZN(
        n20829) );
  OAI22_X1 U12271 ( .A1(n20373), .A2(n25932), .B1(n26219), .B2(n24840), .ZN(
        n20830) );
  OAI22_X1 U12272 ( .A1(n20308), .A2(n25932), .B1(n26218), .B2(n24840), .ZN(
        n20831) );
  OAI22_X1 U12273 ( .A1(n25932), .A2(n28372), .B1(n26192), .B2(n24840), .ZN(
        n22714) );
  OAI22_X1 U12274 ( .A1(n25932), .A2(n28364), .B1(n26193), .B2(n24840), .ZN(
        n22722) );
  OAI22_X1 U12275 ( .A1(n20522), .A2(n25930), .B1(n26221), .B2(n24839), .ZN(
        n20860) );
  OAI22_X1 U12276 ( .A1(n20456), .A2(n25930), .B1(n26220), .B2(n24839), .ZN(
        n20861) );
  OAI22_X1 U12277 ( .A1(n20391), .A2(n25929), .B1(n26219), .B2(n24839), .ZN(
        n20862) );
  OAI22_X1 U12278 ( .A1(n20326), .A2(n25929), .B1(n26218), .B2(n24839), .ZN(
        n20863) );
  OAI22_X1 U12279 ( .A1(n25929), .A2(n28376), .B1(n26192), .B2(n24839), .ZN(
        n22718) );
  OAI22_X1 U12280 ( .A1(n25929), .A2(n28368), .B1(n26193), .B2(n24839), .ZN(
        n22726) );
  OAI22_X1 U12281 ( .A1(n20514), .A2(n25927), .B1(n26251), .B2(n24838), .ZN(
        n20892) );
  OAI22_X1 U12282 ( .A1(n20448), .A2(n25927), .B1(n26250), .B2(n24838), .ZN(
        n20893) );
  OAI22_X1 U12283 ( .A1(n20383), .A2(n25926), .B1(n26249), .B2(n24838), .ZN(
        n20894) );
  OAI22_X1 U12284 ( .A1(n20318), .A2(n25926), .B1(n26248), .B2(n24838), .ZN(
        n20895) );
  OAI22_X1 U12285 ( .A1(n25926), .A2(n28246), .B1(n26252), .B2(n24838), .ZN(
        n22584) );
  OAI22_X1 U12286 ( .A1(n25926), .A2(n28238), .B1(n26253), .B2(n24838), .ZN(
        n22592) );
  OAI22_X1 U12287 ( .A1(n20506), .A2(n25924), .B1(n26221), .B2(n24837), .ZN(
        n20924) );
  OAI22_X1 U12288 ( .A1(n20440), .A2(n25924), .B1(n26220), .B2(n24837), .ZN(
        n20925) );
  OAI22_X1 U12289 ( .A1(n20375), .A2(n25923), .B1(n26219), .B2(n24837), .ZN(
        n20926) );
  OAI22_X1 U12290 ( .A1(n20310), .A2(n25923), .B1(n26218), .B2(n24837), .ZN(
        n20927) );
  OAI22_X1 U12291 ( .A1(n25923), .A2(n28370), .B1(n26192), .B2(n24837), .ZN(
        n22712) );
  OAI22_X1 U12292 ( .A1(n25923), .A2(n28362), .B1(n26193), .B2(n24837), .ZN(
        n22720) );
  OAI22_X1 U12293 ( .A1(n20521), .A2(n25921), .B1(n26221), .B2(n24836), .ZN(
        n20956) );
  OAI22_X1 U12294 ( .A1(n20455), .A2(n25921), .B1(n26220), .B2(n24836), .ZN(
        n20957) );
  OAI22_X1 U12295 ( .A1(n20390), .A2(n25920), .B1(n26219), .B2(n24836), .ZN(
        n20958) );
  OAI22_X1 U12296 ( .A1(n20325), .A2(n25920), .B1(n26218), .B2(n24836), .ZN(
        n20959) );
  OAI22_X1 U12297 ( .A1(n25920), .A2(n28374), .B1(n26192), .B2(n24836), .ZN(
        n22716) );
  OAI22_X1 U12298 ( .A1(n25920), .A2(n28366), .B1(n26193), .B2(n24836), .ZN(
        n22724) );
  OAI22_X1 U12299 ( .A1(n20505), .A2(n25912), .B1(n26221), .B2(n24835), .ZN(
        n21052) );
  OAI22_X1 U12300 ( .A1(n20439), .A2(n25912), .B1(n26220), .B2(n24835), .ZN(
        n21053) );
  OAI22_X1 U12301 ( .A1(n20374), .A2(n25911), .B1(n26219), .B2(n24835), .ZN(
        n21054) );
  OAI22_X1 U12302 ( .A1(n20309), .A2(n25911), .B1(n26218), .B2(n24835), .ZN(
        n21055) );
  OAI22_X1 U12303 ( .A1(n25911), .A2(n28371), .B1(n26192), .B2(n24835), .ZN(
        n22713) );
  OAI22_X1 U12304 ( .A1(n25911), .A2(n28363), .B1(n26193), .B2(n24835), .ZN(
        n22721) );
  OAI22_X1 U12305 ( .A1(n20431), .A2(n25918), .B1(n26220), .B2(n24834), .ZN(
        n20989) );
  OAI22_X1 U12306 ( .A1(n20301), .A2(n25917), .B1(n26218), .B2(n24834), .ZN(
        n20991) );
  OAI22_X1 U12307 ( .A1(n20236), .A2(n25917), .B1(n26217), .B2(n24834), .ZN(
        n20992) );
  OAI22_X1 U12308 ( .A1(n20171), .A2(n25917), .B1(n26216), .B2(n24834), .ZN(
        n20993) );
  OAI22_X1 U12309 ( .A1(n20106), .A2(n25917), .B1(n26215), .B2(n24834), .ZN(
        n20994) );
  OAI22_X1 U12310 ( .A1(n20041), .A2(n25917), .B1(n26214), .B2(n24834), .ZN(
        n20995) );
  INV_X8 U12311 ( .A(n12153), .ZN(n25909) );
  NAND2_X4 U12312 ( .A1(n13093), .A2(n15521), .ZN(n12153) );
endmodule

